module CSRFile(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip,
  input  [11:0] io_rw_addr,
  input  [2:0] io_rw_cmd,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  output  io_csr_stall,
  output  io_csr_xcpt,
  output  io_eret,
  output  io_singleStep,
  output  io_status_debug,
  output [1:0] io_status_prv,
  output  io_status_sd,
  output [30:0] io_status_zero3,
  output  io_status_sd_rv32,
  output [1:0] io_status_zero2,
  output [4:0] io_status_vm,
  output [4:0] io_status_zero1,
  output  io_status_pum,
  output  io_status_mprv,
  output [1:0] io_status_xs,
  output [1:0] io_status_fs,
  output [1:0] io_status_mpp,
  output [1:0] io_status_hpp,
  output  io_status_spp,
  output  io_status_mpie,
  output  io_status_hpie,
  output  io_status_spie,
  output  io_status_upie,
  output  io_status_mie,
  output  io_status_hie,
  output  io_status_sie,
  output  io_status_uie,
  output [6:0] io_ptbr_asid,
  output [37:0] io_ptbr_ppn,
  output [39:0] io_evec,
  input   io_exception,
  input   io_retire,
  input   io_uarch_counters_0,
  input   io_uarch_counters_1,
  input   io_uarch_counters_2,
  input   io_uarch_counters_3,
  input   io_uarch_counters_4,
  input   io_uarch_counters_5,
  input   io_uarch_counters_6,
  input   io_uarch_counters_7,
  input   io_uarch_counters_8,
  input   io_uarch_counters_9,
  input   io_uarch_counters_10,
  input   io_uarch_counters_11,
  input   io_uarch_counters_12,
  input   io_uarch_counters_13,
  input   io_uarch_counters_14,
  input   io_uarch_counters_15,
  input  [63:0] io_cause,
  input  [39:0] io_pc,
  input  [39:0] io_badaddr,
  output  io_fatc,
  output [63:0] io_time,
  output [2:0] io_fcsr_rm,
  input   io_fcsr_flags_valid,
  input  [4:0] io_fcsr_flags_bits,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [63:0] io_rocc_cmd_bits_rs1,
  output [63:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [63:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [39:0] io_rocc_mem_req_bits_addr,
  input  [8:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [63:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [63:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [39:0] io_rocc_mem_resp_bits_addr,
  output [8:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [63:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [63:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  output  io_rocc_status_debug,
  output [1:0] io_rocc_status_prv,
  output  io_rocc_status_sd,
  output [30:0] io_rocc_status_zero3,
  output  io_rocc_status_sd_rv32,
  output [1:0] io_rocc_status_zero2,
  output [4:0] io_rocc_status_vm,
  output [4:0] io_rocc_status_zero1,
  output  io_rocc_status_pum,
  output  io_rocc_status_mprv,
  output [1:0] io_rocc_status_xs,
  output [1:0] io_rocc_status_fs,
  output [1:0] io_rocc_status_mpp,
  output [1:0] io_rocc_status_hpp,
  output  io_rocc_status_spp,
  output  io_rocc_status_mpie,
  output  io_rocc_status_hpie,
  output  io_rocc_status_spie,
  output  io_rocc_status_upie,
  output  io_rocc_status_mie,
  output  io_rocc_status_hie,
  output  io_rocc_status_sie,
  output  io_rocc_status_uie,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input  [1:0] io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [11:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output [1:0] io_rocc_autl_grant_bits_client_xact_id,
  output [2:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception,
  output [11:0] io_rocc_csr_waddr,
  output [63:0] io_rocc_csr_wdata,
  output  io_rocc_csr_wen,
  output  io_rocc_host_id,
  output  io_interrupt,
  output [63:0] io_interrupt_cause,
  output [3:0] io_bp_0_control_tdrtype,
  output [4:0] io_bp_0_control_bpamaskmax,
  output [35:0] io_bp_0_control_reserved,
  output [7:0] io_bp_0_control_bpaction,
  output [3:0] io_bp_0_control_bpmatch,
  output  io_bp_0_control_m,
  output  io_bp_0_control_h,
  output  io_bp_0_control_s,
  output  io_bp_0_control_u,
  output  io_bp_0_control_r,
  output  io_bp_0_control_w,
  output  io_bp_0_control_x,
  output [38:0] io_bp_0_address
);
  wire  T_4992_debug;
  wire [1:0] T_4992_prv;
  wire  T_4992_sd;
  wire [30:0] T_4992_zero3;
  wire  T_4992_sd_rv32;
  wire [1:0] T_4992_zero2;
  wire [4:0] T_4992_vm;
  wire [4:0] T_4992_zero1;
  wire  T_4992_pum;
  wire  T_4992_mprv;
  wire [1:0] T_4992_xs;
  wire [1:0] T_4992_fs;
  wire [1:0] T_4992_mpp;
  wire [1:0] T_4992_hpp;
  wire  T_4992_spp;
  wire  T_4992_mpie;
  wire  T_4992_hpie;
  wire  T_4992_spie;
  wire  T_4992_upie;
  wire  T_4992_mie;
  wire  T_4992_hie;
  wire  T_4992_sie;
  wire  T_4992_uie;
  wire [66:0] T_5017;
  wire  T_5018;
  wire  T_5019;
  wire  T_5020;
  wire  T_5021;
  wire  T_5022;
  wire  T_5023;
  wire  T_5024;
  wire  T_5025;
  wire  T_5026;
  wire [1:0] T_5027;
  wire [1:0] T_5028;
  wire [1:0] T_5029;
  wire [1:0] T_5030;
  wire  T_5031;
  wire  T_5032;
  wire [4:0] T_5033;
  wire [4:0] T_5034;
  wire [1:0] T_5035;
  wire  T_5036;
  wire [30:0] T_5037;
  wire  T_5038;
  wire [1:0] T_5039;
  wire  T_5040;
  wire  reset_mstatus_debug;
  wire [1:0] reset_mstatus_prv;
  wire  reset_mstatus_sd;
  wire [30:0] reset_mstatus_zero3;
  wire  reset_mstatus_sd_rv32;
  wire [1:0] reset_mstatus_zero2;
  wire [4:0] reset_mstatus_vm;
  wire [4:0] reset_mstatus_zero1;
  wire  reset_mstatus_pum;
  wire  reset_mstatus_mprv;
  wire [1:0] reset_mstatus_xs;
  wire [1:0] reset_mstatus_fs;
  wire [1:0] reset_mstatus_mpp;
  wire [1:0] reset_mstatus_hpp;
  wire  reset_mstatus_spp;
  wire  reset_mstatus_mpie;
  wire  reset_mstatus_hpie;
  wire  reset_mstatus_spie;
  wire  reset_mstatus_upie;
  wire  reset_mstatus_mie;
  wire  reset_mstatus_hie;
  wire  reset_mstatus_sie;
  wire  reset_mstatus_uie;
  reg  reg_mstatus_debug;
  reg [31:0] GEN_235;
  reg [1:0] reg_mstatus_prv;
  reg [31:0] GEN_236;
  reg  reg_mstatus_sd;
  reg [31:0] GEN_237;
  reg [30:0] reg_mstatus_zero3;
  reg [31:0] GEN_238;
  reg  reg_mstatus_sd_rv32;
  reg [31:0] GEN_239;
  reg [1:0] reg_mstatus_zero2;
  reg [31:0] GEN_240;
  reg [4:0] reg_mstatus_vm;
  reg [31:0] GEN_241;
  reg [4:0] reg_mstatus_zero1;
  reg [31:0] GEN_242;
  reg  reg_mstatus_pum;
  reg [31:0] GEN_243;
  reg  reg_mstatus_mprv;
  reg [31:0] GEN_244;
  reg [1:0] reg_mstatus_xs;
  reg [31:0] GEN_245;
  reg [1:0] reg_mstatus_fs;
  reg [31:0] GEN_246;
  reg [1:0] reg_mstatus_mpp;
  reg [31:0] GEN_252;
  reg [1:0] reg_mstatus_hpp;
  reg [31:0] GEN_253;
  reg  reg_mstatus_spp;
  reg [31:0] GEN_254;
  reg  reg_mstatus_mpie;
  reg [31:0] GEN_255;
  reg  reg_mstatus_hpie;
  reg [31:0] GEN_256;
  reg  reg_mstatus_spie;
  reg [31:0] GEN_257;
  reg  reg_mstatus_upie;
  reg [31:0] GEN_258;
  reg  reg_mstatus_mie;
  reg [31:0] GEN_259;
  reg  reg_mstatus_hie;
  reg [31:0] GEN_260;
  reg  reg_mstatus_sie;
  reg [31:0] GEN_261;
  reg  reg_mstatus_uie;
  reg [31:0] GEN_262;
  wire [1:0] T_5126_xdebugver;
  wire  T_5126_ndreset;
  wire  T_5126_fullreset;
  wire [11:0] T_5126_hwbpcount;
  wire  T_5126_ebreakm;
  wire  T_5126_ebreakh;
  wire  T_5126_ebreaks;
  wire  T_5126_ebreaku;
  wire  T_5126_zero2;
  wire  T_5126_stopcycle;
  wire  T_5126_stoptime;
  wire [2:0] T_5126_cause;
  wire  T_5126_debugint;
  wire  T_5126_zero1;
  wire  T_5126_halt;
  wire  T_5126_step;
  wire [1:0] T_5126_prv;
  wire [31:0] T_5145;
  wire [1:0] T_5146;
  wire  T_5147;
  wire  T_5148;
  wire  T_5149;
  wire  T_5150;
  wire [2:0] T_5151;
  wire  T_5152;
  wire  T_5153;
  wire  T_5154;
  wire  T_5155;
  wire  T_5156;
  wire  T_5157;
  wire  T_5158;
  wire [11:0] T_5159;
  wire  T_5160;
  wire  T_5161;
  wire [1:0] T_5162;
  wire [1:0] reset_dcsr_xdebugver;
  wire  reset_dcsr_ndreset;
  wire  reset_dcsr_fullreset;
  wire [11:0] reset_dcsr_hwbpcount;
  wire  reset_dcsr_ebreakm;
  wire  reset_dcsr_ebreakh;
  wire  reset_dcsr_ebreaks;
  wire  reset_dcsr_ebreaku;
  wire  reset_dcsr_zero2;
  wire  reset_dcsr_stopcycle;
  wire  reset_dcsr_stoptime;
  wire [2:0] reset_dcsr_cause;
  wire  reset_dcsr_debugint;
  wire  reset_dcsr_zero1;
  wire  reset_dcsr_halt;
  wire  reset_dcsr_step;
  wire [1:0] reset_dcsr_prv;
  reg [1:0] reg_dcsr_xdebugver;
  reg [31:0] GEN_263;
  reg  reg_dcsr_ndreset;
  reg [31:0] GEN_264;
  reg  reg_dcsr_fullreset;
  reg [31:0] GEN_276;
  reg [11:0] reg_dcsr_hwbpcount;
  reg [31:0] GEN_277;
  reg  reg_dcsr_ebreakm;
  reg [31:0] GEN_278;
  reg  reg_dcsr_ebreakh;
  reg [31:0] GEN_279;
  reg  reg_dcsr_ebreaks;
  reg [31:0] GEN_280;
  reg  reg_dcsr_ebreaku;
  reg [31:0] GEN_281;
  reg  reg_dcsr_zero2;
  reg [31:0] GEN_282;
  reg  reg_dcsr_stopcycle;
  reg [31:0] GEN_283;
  reg  reg_dcsr_stoptime;
  reg [31:0] GEN_285;
  reg [2:0] reg_dcsr_cause;
  reg [31:0] GEN_287;
  reg  reg_dcsr_debugint;
  reg [31:0] GEN_288;
  reg  reg_dcsr_zero1;
  reg [31:0] GEN_289;
  reg  reg_dcsr_halt;
  reg [31:0] GEN_291;
  reg  reg_dcsr_step;
  reg [31:0] GEN_293;
  reg [1:0] reg_dcsr_prv;
  reg [31:0] GEN_295;
  wire  T_5228_rocc;
  wire  T_5228_meip;
  wire  T_5228_heip;
  wire  T_5228_seip;
  wire  T_5228_ueip;
  wire  T_5228_mtip;
  wire  T_5228_htip;
  wire  T_5228_stip;
  wire  T_5228_utip;
  wire  T_5228_msip;
  wire  T_5228_hsip;
  wire  T_5228_ssip;
  wire  T_5228_usip;
  wire [12:0] T_5243;
  wire  T_5244;
  wire  T_5245;
  wire  T_5246;
  wire  T_5247;
  wire  T_5248;
  wire  T_5249;
  wire  T_5250;
  wire  T_5251;
  wire  T_5252;
  wire  T_5253;
  wire  T_5254;
  wire  T_5255;
  wire  T_5256;
  wire  T_5257_rocc;
  wire  T_5257_meip;
  wire  T_5257_heip;
  wire  T_5257_seip;
  wire  T_5257_ueip;
  wire  T_5257_mtip;
  wire  T_5257_htip;
  wire  T_5257_stip;
  wire  T_5257_utip;
  wire  T_5257_msip;
  wire  T_5257_hsip;
  wire  T_5257_ssip;
  wire  T_5257_usip;
  wire  T_5278_rocc;
  wire  T_5278_meip;
  wire  T_5278_heip;
  wire  T_5278_seip;
  wire  T_5278_ueip;
  wire  T_5278_mtip;
  wire  T_5278_htip;
  wire  T_5278_stip;
  wire  T_5278_utip;
  wire  T_5278_msip;
  wire  T_5278_hsip;
  wire  T_5278_ssip;
  wire  T_5278_usip;
  wire [1:0] T_5295;
  wire [2:0] T_5296;
  wire [1:0] T_5297;
  wire [2:0] T_5298;
  wire [5:0] T_5299;
  wire [1:0] T_5300;
  wire [2:0] T_5301;
  wire [1:0] T_5302;
  wire [1:0] T_5303;
  wire [3:0] T_5304;
  wire [6:0] T_5305;
  wire [12:0] supported_interrupts;
  wire [1:0] T_5306;
  wire [2:0] T_5307;
  wire [1:0] T_5308;
  wire [2:0] T_5309;
  wire [5:0] T_5310;
  wire [1:0] T_5311;
  wire [2:0] T_5312;
  wire [1:0] T_5313;
  wire [1:0] T_5314;
  wire [3:0] T_5315;
  wire [6:0] T_5316;
  wire [12:0] delegable_interrupts;
  wire  exception;
  reg  reg_debug;
  reg [31:0] GEN_297;
  reg [39:0] reg_dpc;
  reg [63:0] GEN_299;
  reg [63:0] reg_dscratch;
  reg [63:0] GEN_301;
  reg  reg_singleStepped;
  reg [31:0] GEN_302;
  wire  T_5322;
  wire  GEN_27;
  wire  T_5325;
  wire  GEN_28;
  wire  T_5336;
  wire  T_5338;
  wire  T_5339;
  wire  T_5340;
  wire  T_5342;
  reg  reg_tdrselect_tdrmode;
  reg [31:0] GEN_303;
  reg [61:0] reg_tdrselect_reserved;
  reg [63:0] GEN_304;
  reg  reg_tdrselect_tdrindex;
  reg [31:0] GEN_305;
  reg [3:0] reg_bp_0_control_tdrtype;
  reg [31:0] GEN_306;
  reg [4:0] reg_bp_0_control_bpamaskmax;
  reg [31:0] GEN_307;
  reg [35:0] reg_bp_0_control_reserved;
  reg [63:0] GEN_308;
  reg [7:0] reg_bp_0_control_bpaction;
  reg [31:0] GEN_309;
  reg [3:0] reg_bp_0_control_bpmatch;
  reg [31:0] GEN_310;
  reg  reg_bp_0_control_m;
  reg [31:0] GEN_311;
  reg  reg_bp_0_control_h;
  reg [31:0] GEN_312;
  reg  reg_bp_0_control_s;
  reg [31:0] GEN_313;
  reg  reg_bp_0_control_u;
  reg [31:0] GEN_314;
  reg  reg_bp_0_control_r;
  reg [31:0] GEN_315;
  reg  reg_bp_0_control_w;
  reg [31:0] GEN_316;
  reg  reg_bp_0_control_x;
  reg [31:0] GEN_317;
  reg [38:0] reg_bp_0_address;
  reg [63:0] GEN_318;
  reg [3:0] reg_bp_1_control_tdrtype;
  reg [31:0] GEN_319;
  reg [4:0] reg_bp_1_control_bpamaskmax;
  reg [31:0] GEN_320;
  reg [35:0] reg_bp_1_control_reserved;
  reg [63:0] GEN_321;
  reg [7:0] reg_bp_1_control_bpaction;
  reg [31:0] GEN_322;
  reg [3:0] reg_bp_1_control_bpmatch;
  reg [31:0] GEN_323;
  reg  reg_bp_1_control_m;
  reg [31:0] GEN_324;
  reg  reg_bp_1_control_h;
  reg [31:0] GEN_325;
  reg  reg_bp_1_control_s;
  reg [31:0] GEN_326;
  reg  reg_bp_1_control_u;
  reg [31:0] GEN_328;
  reg  reg_bp_1_control_r;
  reg [31:0] GEN_329;
  reg  reg_bp_1_control_w;
  reg [31:0] GEN_331;
  reg  reg_bp_1_control_x;
  reg [31:0] GEN_332;
  reg [38:0] reg_bp_1_address;
  reg [63:0] GEN_333;
  reg [63:0] reg_mie;
  reg [63:0] GEN_334;
  reg [63:0] reg_mideleg;
  reg [63:0] GEN_335;
  reg [63:0] reg_medeleg;
  reg [63:0] GEN_337;
  reg  reg_mip_rocc;
  reg [31:0] GEN_338;
  reg  reg_mip_meip;
  reg [31:0] GEN_340;
  reg  reg_mip_heip;
  reg [31:0] GEN_341;
  reg  reg_mip_seip;
  reg [31:0] GEN_343;
  reg  reg_mip_ueip;
  reg [31:0] GEN_344;
  reg  reg_mip_mtip;
  reg [31:0] GEN_346;
  reg  reg_mip_htip;
  reg [31:0] GEN_347;
  reg  reg_mip_stip;
  reg [31:0] GEN_349;
  reg  reg_mip_utip;
  reg [31:0] GEN_350;
  reg  reg_mip_msip;
  reg [31:0] GEN_352;
  reg  reg_mip_hsip;
  reg [31:0] GEN_353;
  reg  reg_mip_ssip;
  reg [31:0] GEN_355;
  reg  reg_mip_usip;
  reg [31:0] GEN_356;
  reg [39:0] reg_mepc;
  reg [63:0] GEN_357;
  reg [63:0] reg_mcause;
  reg [63:0] GEN_358;
  reg [39:0] reg_mbadaddr;
  reg [63:0] GEN_359;
  reg [63:0] reg_mscratch;
  reg [63:0] GEN_360;
  reg [31:0] reg_mtvec;
  reg [31:0] GEN_361;
  reg [39:0] reg_sepc;
  reg [63:0] GEN_362;
  reg [63:0] reg_scause;
  reg [63:0] GEN_363;
  reg [39:0] reg_sbadaddr;
  reg [63:0] GEN_364;
  reg [63:0] reg_sscratch;
  reg [63:0] GEN_365;
  reg [38:0] reg_stvec;
  reg [63:0] GEN_366;
  reg [6:0] reg_sptbr_asid;
  reg [31:0] GEN_367;
  reg [37:0] reg_sptbr_ppn;
  reg [63:0] GEN_368;
  reg  reg_wfi;
  reg [31:0] GEN_369;
  reg [5:0] T_5544;
  reg [31:0] GEN_370;
  wire [6:0] GEN_595;
  wire [7:0] T_5548;
  wire [6:0] T_5549;
  wire [5:0] T_5550;
  wire [5:0] GEN_29;
  reg [57:0] T_5552;
  reg [63:0] GEN_371;
  wire  T_5553;
  wire  T_5554;
  wire [57:0] GEN_596;
  wire [58:0] T_5556;
  wire [57:0] T_5557;
  wire [57:0] GEN_30;
  reg [5:0] T_5560;
  reg [31:0] GEN_372;
  wire [6:0] GEN_597;
  wire [7:0] T_5564;
  wire [6:0] T_5565;
  wire [5:0] T_5566;
  wire [5:0] GEN_31;
  reg [57:0] T_5568;
  reg [63:0] GEN_373;
  wire  T_5569;
  wire  T_5570;
  wire [58:0] T_5572;
  wire [57:0] T_5573;
  wire [57:0] GEN_32;
  reg [5:0] T_5576;
  reg [31:0] GEN_374;
  wire [6:0] GEN_599;
  wire [7:0] T_5580;
  wire [6:0] T_5581;
  wire [5:0] T_5582;
  wire [5:0] GEN_33;
  reg [57:0] T_5584;
  reg [63:0] GEN_375;
  wire  T_5585;
  wire  T_5586;
  wire [58:0] T_5588;
  wire [57:0] T_5589;
  wire [57:0] GEN_34;
  reg [5:0] T_5592;
  reg [31:0] GEN_376;
  wire [6:0] GEN_601;
  wire [7:0] T_5596;
  wire [6:0] T_5597;
  wire [5:0] T_5598;
  wire [5:0] GEN_35;
  reg [57:0] T_5600;
  reg [63:0] GEN_377;
  wire  T_5601;
  wire  T_5602;
  wire [58:0] T_5604;
  wire [57:0] T_5605;
  wire [57:0] GEN_36;
  reg [5:0] T_5608;
  reg [31:0] GEN_378;
  wire [6:0] GEN_603;
  wire [7:0] T_5612;
  wire [6:0] T_5613;
  wire [5:0] T_5614;
  wire [5:0] GEN_37;
  reg [57:0] T_5616;
  reg [63:0] GEN_379;
  wire  T_5617;
  wire  T_5618;
  wire [58:0] T_5620;
  wire [57:0] T_5621;
  wire [57:0] GEN_38;
  reg [5:0] T_5624;
  reg [31:0] GEN_380;
  wire [6:0] GEN_605;
  wire [7:0] T_5628;
  wire [6:0] T_5629;
  wire [5:0] T_5630;
  wire [5:0] GEN_39;
  reg [57:0] T_5632;
  reg [63:0] GEN_382;
  wire  T_5633;
  wire  T_5634;
  wire [58:0] T_5636;
  wire [57:0] T_5637;
  wire [57:0] GEN_40;
  reg [5:0] T_5640;
  reg [31:0] GEN_383;
  wire [6:0] GEN_607;
  wire [7:0] T_5644;
  wire [6:0] T_5645;
  wire [5:0] T_5646;
  wire [5:0] GEN_41;
  reg [57:0] T_5648;
  reg [63:0] GEN_385;
  wire  T_5649;
  wire  T_5650;
  wire [58:0] T_5652;
  wire [57:0] T_5653;
  wire [57:0] GEN_42;
  reg [5:0] T_5656;
  reg [31:0] GEN_386;
  wire [6:0] GEN_609;
  wire [7:0] T_5660;
  wire [6:0] T_5661;
  wire [5:0] T_5662;
  wire [5:0] GEN_43;
  reg [57:0] T_5664;
  reg [63:0] GEN_387;
  wire  T_5665;
  wire  T_5666;
  wire [58:0] T_5668;
  wire [57:0] T_5669;
  wire [57:0] GEN_44;
  reg [5:0] T_5672;
  reg [31:0] GEN_388;
  wire [6:0] GEN_611;
  wire [7:0] T_5676;
  wire [6:0] T_5677;
  wire [5:0] T_5678;
  wire [5:0] GEN_45;
  reg [57:0] T_5680;
  reg [63:0] GEN_389;
  wire  T_5681;
  wire  T_5682;
  wire [58:0] T_5684;
  wire [57:0] T_5685;
  wire [57:0] GEN_46;
  reg [5:0] T_5688;
  reg [31:0] GEN_391;
  wire [6:0] GEN_613;
  wire [7:0] T_5692;
  wire [6:0] T_5693;
  wire [5:0] T_5694;
  wire [5:0] GEN_47;
  reg [57:0] T_5696;
  reg [63:0] GEN_392;
  wire  T_5697;
  wire  T_5698;
  wire [58:0] T_5700;
  wire [57:0] T_5701;
  wire [57:0] GEN_48;
  reg [5:0] T_5704;
  reg [31:0] GEN_394;
  wire [6:0] GEN_615;
  wire [7:0] T_5708;
  wire [6:0] T_5709;
  wire [5:0] T_5710;
  wire [5:0] GEN_49;
  reg [57:0] T_5712;
  reg [63:0] GEN_395;
  wire  T_5713;
  wire  T_5714;
  wire [58:0] T_5716;
  wire [57:0] T_5717;
  wire [57:0] GEN_50;
  reg [5:0] T_5720;
  reg [31:0] GEN_397;
  wire [6:0] GEN_617;
  wire [7:0] T_5724;
  wire [6:0] T_5725;
  wire [5:0] T_5726;
  wire [5:0] GEN_51;
  reg [57:0] T_5728;
  reg [63:0] GEN_398;
  wire  T_5729;
  wire  T_5730;
  wire [58:0] T_5732;
  wire [57:0] T_5733;
  wire [57:0] GEN_52;
  reg [5:0] T_5736;
  reg [31:0] GEN_400;
  wire [6:0] GEN_619;
  wire [7:0] T_5740;
  wire [6:0] T_5741;
  wire [5:0] T_5742;
  wire [5:0] GEN_53;
  reg [57:0] T_5744;
  reg [63:0] GEN_401;
  wire  T_5745;
  wire  T_5746;
  wire [58:0] T_5748;
  wire [57:0] T_5749;
  wire [57:0] GEN_54;
  reg [5:0] T_5752;
  reg [31:0] GEN_403;
  wire [6:0] GEN_621;
  wire [7:0] T_5756;
  wire [6:0] T_5757;
  wire [5:0] T_5758;
  wire [5:0] GEN_55;
  reg [57:0] T_5760;
  reg [63:0] GEN_404;
  wire  T_5761;
  wire  T_5762;
  wire [58:0] T_5764;
  wire [57:0] T_5765;
  wire [57:0] GEN_56;
  reg [5:0] T_5768;
  reg [31:0] GEN_405;
  wire [6:0] GEN_623;
  wire [7:0] T_5772;
  wire [6:0] T_5773;
  wire [5:0] T_5774;
  wire [5:0] GEN_57;
  reg [57:0] T_5776;
  reg [63:0] GEN_407;
  wire  T_5777;
  wire  T_5778;
  wire [58:0] T_5780;
  wire [57:0] T_5781;
  wire [57:0] GEN_58;
  reg [5:0] T_5784;
  reg [31:0] GEN_408;
  wire [6:0] GEN_625;
  wire [7:0] T_5788;
  wire [6:0] T_5789;
  wire [5:0] T_5790;
  wire [5:0] GEN_59;
  reg [57:0] T_5792;
  reg [63:0] GEN_409;
  wire  T_5793;
  wire  T_5794;
  wire [58:0] T_5796;
  wire [57:0] T_5797;
  wire [57:0] GEN_60;
  reg [4:0] reg_fflags;
  reg [31:0] GEN_410;
  reg [2:0] reg_frm;
  reg [31:0] GEN_411;
  reg [5:0] T_5802;
  reg [31:0] GEN_412;
  wire [6:0] GEN_627;
  wire [7:0] T_5806;
  wire [6:0] T_5807;
  wire [5:0] T_5808;
  wire [5:0] GEN_61;
  reg [57:0] T_5810;
  reg [63:0] GEN_413;
  wire  T_5811;
  wire  T_5812;
  wire [58:0] T_5814;
  wire [57:0] T_5815;
  wire [57:0] GEN_62;
  wire [63:0] T_5816;
  reg [5:0] T_5819;
  reg [31:0] GEN_414;
  wire [6:0] GEN_629;
  wire [7:0] T_5823;
  wire [6:0] T_5824;
  wire [5:0] T_5825;
  reg [57:0] T_5827;
  reg [63:0] GEN_415;
  wire  T_5828;
  wire [58:0] T_5831;
  wire [57:0] T_5832;
  wire [57:0] GEN_64;
  wire [63:0] reg_cycle;
  wire  mip_rocc;
  wire  mip_meip;
  wire  mip_heip;
  wire  mip_seip;
  wire  mip_ueip;
  wire  mip_mtip;
  wire  mip_htip;
  wire  mip_stip;
  wire  mip_utip;
  wire  mip_msip;
  wire  mip_hsip;
  wire  mip_ssip;
  wire  mip_usip;
  wire [1:0] T_5846;
  wire [2:0] T_5847;
  wire [1:0] T_5848;
  wire [2:0] T_5849;
  wire [5:0] T_5850;
  wire [1:0] T_5851;
  wire [2:0] T_5852;
  wire [1:0] T_5853;
  wire [1:0] T_5854;
  wire [3:0] T_5855;
  wire [6:0] T_5856;
  wire [12:0] T_5857;
  wire [12:0] read_mip;
  wire [63:0] GEN_631;
  wire [63:0] pending_interrupts;
  wire  T_5859;
  wire  T_5861;
  wire  T_5863;
  wire  T_5864;
  wire  T_5865;
  wire  T_5866;
  wire [63:0] T_5867;
  wire [63:0] T_5868;
  wire [63:0] m_interrupts;
  wire [1:0] GEN_632;
  wire  T_5873;
  wire  T_5875;
  wire  T_5876;
  wire  T_5877;
  wire  T_5878;
  wire [63:0] T_5879;
  wire [63:0] s_interrupts;
  wire [63:0] all_interrupts;
  wire  T_5882;
  wire  T_5883;
  wire  T_5884;
  wire  T_5885;
  wire  T_5886;
  wire  T_5887;
  wire  T_5888;
  wire  T_5889;
  wire  T_5890;
  wire  T_5891;
  wire  T_5892;
  wire  T_5893;
  wire  T_5894;
  wire  T_5895;
  wire  T_5896;
  wire  T_5897;
  wire  T_5898;
  wire  T_5899;
  wire  T_5900;
  wire  T_5901;
  wire  T_5902;
  wire  T_5903;
  wire  T_5904;
  wire  T_5905;
  wire  T_5906;
  wire  T_5907;
  wire  T_5908;
  wire  T_5909;
  wire  T_5910;
  wire  T_5911;
  wire  T_5912;
  wire  T_5913;
  wire  T_5914;
  wire  T_5915;
  wire  T_5916;
  wire  T_5917;
  wire  T_5918;
  wire  T_5919;
  wire  T_5920;
  wire  T_5921;
  wire  T_5922;
  wire  T_5923;
  wire  T_5924;
  wire  T_5925;
  wire  T_5926;
  wire  T_5927;
  wire  T_5928;
  wire  T_5929;
  wire  T_5930;
  wire  T_5931;
  wire  T_5932;
  wire  T_5933;
  wire  T_5934;
  wire  T_5935;
  wire  T_5936;
  wire  T_5937;
  wire  T_5938;
  wire  T_5939;
  wire  T_5940;
  wire  T_5941;
  wire  T_5942;
  wire  T_5943;
  wire  T_5944;
  wire [5:0] T_6010;
  wire [5:0] T_6011;
  wire [5:0] T_6012;
  wire [5:0] T_6013;
  wire [5:0] T_6014;
  wire [5:0] T_6015;
  wire [5:0] T_6016;
  wire [5:0] T_6017;
  wire [5:0] T_6018;
  wire [5:0] T_6019;
  wire [5:0] T_6020;
  wire [5:0] T_6021;
  wire [5:0] T_6022;
  wire [5:0] T_6023;
  wire [5:0] T_6024;
  wire [5:0] T_6025;
  wire [5:0] T_6026;
  wire [5:0] T_6027;
  wire [5:0] T_6028;
  wire [5:0] T_6029;
  wire [5:0] T_6030;
  wire [5:0] T_6031;
  wire [5:0] T_6032;
  wire [5:0] T_6033;
  wire [5:0] T_6034;
  wire [5:0] T_6035;
  wire [5:0] T_6036;
  wire [5:0] T_6037;
  wire [5:0] T_6038;
  wire [5:0] T_6039;
  wire [5:0] T_6040;
  wire [5:0] T_6041;
  wire [5:0] T_6042;
  wire [5:0] T_6043;
  wire [5:0] T_6044;
  wire [5:0] T_6045;
  wire [5:0] T_6046;
  wire [5:0] T_6047;
  wire [5:0] T_6048;
  wire [5:0] T_6049;
  wire [5:0] T_6050;
  wire [5:0] T_6051;
  wire [5:0] T_6052;
  wire [5:0] T_6053;
  wire [5:0] T_6054;
  wire [5:0] T_6055;
  wire [5:0] T_6056;
  wire [5:0] T_6057;
  wire [5:0] T_6058;
  wire [5:0] T_6059;
  wire [5:0] T_6060;
  wire [5:0] T_6061;
  wire [5:0] T_6062;
  wire [5:0] T_6063;
  wire [5:0] T_6064;
  wire [5:0] T_6065;
  wire [5:0] T_6066;
  wire [5:0] T_6067;
  wire [5:0] T_6068;
  wire [5:0] T_6069;
  wire [5:0] T_6070;
  wire [5:0] T_6071;
  wire [5:0] T_6072;
  wire [63:0] GEN_634;
  wire [64:0] T_6073;
  wire [63:0] interruptCause;
  wire [63:0] GEN_635;
  wire  T_6075;
  wire  T_6078;
  wire  T_6079;
  wire  T_6084;
  wire  GEN_65;
  wire [63:0] GEN_66;
  wire  system_insn;
  wire  T_6087;
  wire  T_6089;
  wire  cpu_ren;
  wire [1:0] T_6090;
  wire [1:0] T_6091;
  wire [2:0] T_6092;
  wire [4:0] T_6093;
  wire [1:0] T_6094;
  wire [2:0] T_6095;
  wire [3:0] T_6096;
  wire [4:0] T_6097;
  wire [7:0] T_6098;
  wire [12:0] T_6099;
  wire [2:0] T_6100;
  wire [4:0] T_6101;
  wire [9:0] T_6102;
  wire [10:0] T_6103;
  wire [15:0] T_6104;
  wire [31:0] T_6105;
  wire [33:0] T_6106;
  wire [2:0] T_6107;
  wire [3:0] T_6108;
  wire [37:0] T_6109;
  wire [53:0] T_6110;
  wire [66:0] T_6111;
  wire [63:0] read_mstatus;
  wire [62:0] T_6112;
  wire [63:0] T_6113;
  wire  GEN_0;
  wire  GEN_67;
  wire  GEN_1;
  wire  GEN_68;
  wire [1:0] T_6128;
  wire  GEN_2;
  wire  GEN_69;
  wire [2:0] T_6129;
  wire  GEN_3;
  wire  GEN_70;
  wire  GEN_4;
  wire  GEN_71;
  wire [1:0] T_6130;
  wire  GEN_5;
  wire  GEN_72;
  wire [2:0] T_6131;
  wire [5:0] T_6132;
  wire [7:0] GEN_6;
  wire [7:0] GEN_73;
  wire [3:0] GEN_7;
  wire [3:0] GEN_74;
  wire [11:0] T_6133;
  wire  GEN_8;
  wire  GEN_75;
  wire [12:0] T_6134;
  wire [3:0] GEN_9;
  wire [3:0] GEN_76;
  wire [4:0] GEN_10;
  wire [4:0] GEN_77;
  wire [8:0] T_6135;
  wire [35:0] GEN_11;
  wire [35:0] GEN_78;
  wire [44:0] T_6136;
  wire [57:0] T_6137;
  wire [63:0] T_6138;
  wire  T_6161;
  wire [23:0] GEN_636;
  wire [24:0] T_6163;
  wire [23:0] T_6164;
  wire [63:0] T_6165;
  wire  T_6166;
  wire [23:0] GEN_637;
  wire [24:0] T_6168;
  wire [23:0] T_6169;
  wire [63:0] T_6170;
  wire [2:0] T_6171;
  wire [1:0] T_6172;
  wire [4:0] T_6173;
  wire [3:0] T_6174;
  wire [1:0] T_6175;
  wire [5:0] T_6176;
  wire [10:0] T_6177;
  wire [1:0] T_6178;
  wire [1:0] T_6179;
  wire [3:0] T_6180;
  wire [12:0] T_6181;
  wire [2:0] T_6182;
  wire [3:0] T_6183;
  wire [16:0] T_6184;
  wire [20:0] T_6185;
  wire [31:0] T_6186;
  wire [63:0] T_6187;
  wire [63:0] T_6188;
  wire  T_6189_debug;
  wire [1:0] T_6189_prv;
  wire  T_6189_sd;
  wire [30:0] T_6189_zero3;
  wire  T_6189_sd_rv32;
  wire [1:0] T_6189_zero2;
  wire [4:0] T_6189_vm;
  wire [4:0] T_6189_zero1;
  wire  T_6189_pum;
  wire  T_6189_mprv;
  wire [1:0] T_6189_xs;
  wire [1:0] T_6189_fs;
  wire [1:0] T_6189_mpp;
  wire [1:0] T_6189_hpp;
  wire  T_6189_spp;
  wire  T_6189_mpie;
  wire  T_6189_hpie;
  wire  T_6189_spie;
  wire  T_6189_upie;
  wire  T_6189_mie;
  wire  T_6189_hie;
  wire  T_6189_sie;
  wire  T_6189_uie;
  wire [1:0] T_6221;
  wire [1:0] T_6222;
  wire [2:0] T_6223;
  wire [4:0] T_6224;
  wire [1:0] T_6225;
  wire [2:0] T_6226;
  wire [3:0] T_6227;
  wire [4:0] T_6228;
  wire [7:0] T_6229;
  wire [12:0] T_6230;
  wire [2:0] T_6231;
  wire [4:0] T_6232;
  wire [9:0] T_6233;
  wire [10:0] T_6234;
  wire [15:0] T_6235;
  wire [31:0] T_6236;
  wire [33:0] T_6237;
  wire [2:0] T_6238;
  wire [3:0] T_6239;
  wire [37:0] T_6240;
  wire [53:0] T_6241;
  wire [66:0] T_6242;
  wire [63:0] T_6243;
  wire  T_6244;
  wire [23:0] GEN_639;
  wire [24:0] T_6246;
  wire [23:0] T_6247;
  wire [63:0] T_6248;
  wire [44:0] T_6249;
  wire  T_6250;
  wire [23:0] GEN_640;
  wire [24:0] T_6252;
  wire [23:0] T_6253;
  wire [63:0] T_6254;
  wire  T_6255;
  wire [24:0] GEN_641;
  wire [25:0] T_6257;
  wire [24:0] T_6258;
  wire [63:0] T_6259;
  wire [11:0] GEN_642;
  wire  T_6265;
  wire [11:0] GEN_643;
  wire  T_6267;
  wire [11:0] GEN_644;
  wire  T_6269;
  wire  T_6271;
  wire  T_6273;
  wire  T_6275;
  wire  T_6277;
  wire  T_6279;
  wire [11:0] GEN_645;
  wire  T_6281;
  wire [11:0] GEN_646;
  wire  T_6283;
  wire [11:0] GEN_647;
  wire  T_6285;
  wire [11:0] GEN_648;
  wire  T_6287;
  wire  T_6289;
  wire [11:0] GEN_649;
  wire  T_6291;
  wire [11:0] GEN_650;
  wire  T_6293;
  wire [11:0] GEN_651;
  wire  T_6295;
  wire [11:0] GEN_652;
  wire  T_6297;
  wire [11:0] GEN_653;
  wire  T_6299;
  wire [11:0] GEN_654;
  wire  T_6301;
  wire [11:0] GEN_655;
  wire  T_6303;
  wire [11:0] GEN_656;
  wire  T_6305;
  wire [11:0] GEN_657;
  wire  T_6307;
  wire [11:0] GEN_658;
  wire  T_6309;
  wire  T_6311;
  wire [11:0] GEN_659;
  wire  T_6313;
  wire [11:0] GEN_660;
  wire  T_6315;
  wire [11:0] GEN_661;
  wire  T_6317;
  wire [11:0] GEN_662;
  wire  T_6319;
  wire [11:0] GEN_663;
  wire  T_6321;
  wire [11:0] GEN_664;
  wire  T_6323;
  wire [11:0] GEN_665;
  wire  T_6325;
  wire [11:0] GEN_666;
  wire  T_6327;
  wire [11:0] GEN_667;
  wire  T_6329;
  wire [11:0] GEN_668;
  wire  T_6331;
  wire [11:0] GEN_669;
  wire  T_6333;
  wire [11:0] GEN_670;
  wire  T_6335;
  wire [11:0] GEN_671;
  wire  T_6337;
  wire [11:0] GEN_672;
  wire  T_6339;
  wire [11:0] GEN_673;
  wire  T_6341;
  wire [11:0] GEN_674;
  wire  T_6343;
  wire  T_6344;
  wire  T_6345;
  wire  T_6346;
  wire  T_6347;
  wire  T_6348;
  wire  T_6349;
  wire  T_6350;
  wire  T_6351;
  wire  T_6352;
  wire  T_6353;
  wire  T_6354;
  wire  T_6355;
  wire  T_6356;
  wire  T_6357;
  wire  T_6358;
  wire  T_6359;
  wire  T_6360;
  wire  T_6361;
  wire  T_6362;
  wire  T_6363;
  wire  T_6364;
  wire  T_6365;
  wire  T_6366;
  wire  T_6367;
  wire  T_6368;
  wire  T_6369;
  wire  T_6370;
  wire  T_6371;
  wire  T_6372;
  wire  T_6373;
  wire  T_6374;
  wire  T_6375;
  wire  T_6376;
  wire  T_6377;
  wire  T_6378;
  wire  T_6379;
  wire  T_6380;
  wire  T_6381;
  wire  addr_valid;
  wire  T_6383;
  wire [1:0] T_6384;
  wire [1:0] T_6385;
  wire [1:0] GEN_675;
  wire  T_6387;
  wire [1:0] T_6388;
  wire [2:0] csr_addr_priv;
  wire [2:0] T_6389;
  wire  priv_sufficient;
  wire [1:0] T_6390;
  wire [1:0] T_6391;
  wire  read_only;
  wire  T_6393;
  wire  T_6394;
  wire  cpu_wen;
  wire  T_6396;
  wire  wen;
  wire  T_6397;
  wire  T_6398;
  wire  T_6399;
  wire [63:0] T_6401;
  wire  T_6402;
  wire [63:0] T_6404;
  wire [63:0] T_6405;
  wire [63:0] T_6408;
  wire [63:0] T_6409;
  wire [63:0] wdata;
  wire  do_system_insn;
  wire [2:0] T_6411;
  wire [7:0] GEN_677;
  wire [7:0] opcode;
  wire  T_6412;
  wire  insn_call;
  wire  T_6413;
  wire  insn_break;
  wire  T_6414;
  wire  insn_ret;
  wire  T_6415;
  wire  insn_sfence_vm;
  wire  T_6416;
  wire  insn_wfi;
  wire  T_6417;
  wire  T_6419;
  wire  T_6421;
  wire  T_6422;
  wire  T_6429;
  wire  T_6430;
  wire  T_6433;
  wire  T_6434;
  wire  T_6435;
  wire  T_6436;
  wire  GEN_79;
  wire [12:0] GEN_679;
  wire  T_6439;
  wire  GEN_80;
  wire  T_6442;
  wire [3:0] GEN_680;
  wire [4:0] T_6444;
  wire [3:0] T_6445;
  wire [1:0] T_6448;
  wire [3:0] T_6449;
  wire [63:0] cause;
  wire [5:0] cause_lsbs;
  wire  T_6450;
  wire [5:0] GEN_681;
  wire  T_6452;
  wire  causeIsDebugInt;
  wire [63:0] GEN_682;
  wire  T_6454;
  wire [1:0] T_6455;
  wire [1:0] T_6456;
  wire [3:0] T_6457;
  wire [3:0] T_6458;
  wire  T_6459;
  wire  causeIsDebugBreak;
  wire  T_6461;
  wire  T_6462;
  wire  T_6463;
  wire [63:0] T_6469;
  wire  T_6470;
  wire [63:0] T_6471;
  wire  T_6472;
  wire  T_6473;
  wire  delegate;
  wire [11:0] debugTVec;
  wire [39:0] T_6477;
  wire [39:0] T_6478;
  wire [39:0] tvec;
  wire  T_6480;
  wire  T_6482;
  wire [39:0] T_6484;
  wire [39:0] epc;
  wire [39:0] T_6485;
  wire  T_6488;
  wire [1:0] T_6489;
  wire  T_6491;
  wire [1:0] T_6492;
  wire  T_6494;
  wire  T_6495;
  wire [39:0] T_6496;
  wire [39:0] GEN_685;
  wire [39:0] T_6498;
  wire [39:0] T_6499;
  wire [63:0] T_6500;
  wire  T_6501;
  wire [1:0] T_6506;
  wire [2:0] T_6507;
  wire  GEN_81;
  wire [39:0] GEN_82;
  wire [2:0] GEN_83;
  wire [1:0] GEN_84;
  wire  T_6509;
  wire  T_6510;
  wire [39:0] GEN_85;
  wire [63:0] GEN_86;
  wire [39:0] GEN_87;
  wire  GEN_88;
  wire [1:0] GEN_89;
  wire  GEN_90;
  wire [1:0] GEN_91;
  wire  T_6516;
  wire  T_6517;
  wire [39:0] GEN_92;
  wire [63:0] GEN_93;
  wire [39:0] GEN_94;
  wire  GEN_95;
  wire [1:0] GEN_96;
  wire  GEN_97;
  wire [1:0] GEN_98;
  wire  GEN_99;
  wire [39:0] GEN_100;
  wire [2:0] GEN_101;
  wire [1:0] GEN_102;
  wire [39:0] GEN_103;
  wire [63:0] GEN_104;
  wire [39:0] GEN_105;
  wire  GEN_106;
  wire [1:0] GEN_107;
  wire  GEN_108;
  wire [1:0] GEN_109;
  wire [39:0] GEN_110;
  wire [63:0] GEN_111;
  wire [39:0] GEN_112;
  wire  GEN_113;
  wire [1:0] GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire [1:0] GEN_119;
  wire [1:0] GEN_120;
  wire  T_6529;
  wire  T_6530;
  wire [1:0] GEN_121;
  wire  GEN_122;
  wire  T_6535;
  wire  T_6536;
  wire  T_6537;
  wire  GEN_123;
  wire  T_6539;
  wire  T_6542;
  wire  T_6543;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire [1:0] GEN_128;
  wire [1:0] GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire [1:0] GEN_132;
  wire [1:0] GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire [1:0] GEN_137;
  wire [1:0] T_6548;
  wire [1:0] GEN_686;
  wire [2:0] T_6549;
  wire [1:0] T_6550;
  wire [2:0] T_6551;
  wire [2:0] GEN_687;
  wire [3:0] T_6552;
  wire [2:0] T_6553;
  wire [2:0] GEN_688;
  wire  T_6555;
  wire  T_6556;
  wire  T_6558;
  wire [63:0] T_6560;
  wire [63:0] T_6562;
  wire [38:0] GEN_12;
  wire [38:0] GEN_138;
  wire [38:0] T_6564;
  wire [63:0] T_6572;
  wire [63:0] T_6574;
  wire [63:0] T_6584;
  wire [63:0] T_6586;
  wire [31:0] T_6588;
  wire [12:0] T_6590;
  wire [63:0] T_6592;
  wire [63:0] T_6594;
  wire [63:0] T_6596;
  wire [63:0] T_6598;
  wire [63:0] T_6600;
  wire [63:0] T_6602;
  wire [63:0] T_6604;
  wire  T_6606;
  wire [31:0] T_6608;
  wire [39:0] T_6610;
  wire [63:0] T_6612;
  wire [63:0] T_6614;
  wire [63:0] T_6616;
  wire [63:0] T_6618;
  wire [63:0] T_6620;
  wire [63:0] T_6622;
  wire [63:0] T_6624;
  wire [44:0] T_6626;
  wire [63:0] T_6628;
  wire [63:0] T_6630;
  wire [63:0] T_6640;
  wire [63:0] GEN_689;
  wire [63:0] T_6641;
  wire [63:0] T_6642;
  wire [63:0] T_6643;
  wire [63:0] T_6644;
  wire [63:0] T_6645;
  wire [63:0] T_6646;
  wire [63:0] T_6647;
  wire [63:0] T_6648;
  wire [63:0] T_6649;
  wire [63:0] T_6650;
  wire [63:0] T_6651;
  wire [63:0] T_6652;
  wire [63:0] GEN_697;
  wire [63:0] T_6653;
  wire [63:0] GEN_698;
  wire [63:0] T_6654;
  wire [63:0] T_6655;
  wire [63:0] T_6656;
  wire [63:0] T_6657;
  wire [63:0] T_6658;
  wire [63:0] T_6659;
  wire [63:0] T_6660;
  wire [63:0] T_6661;
  wire [63:0] GEN_699;
  wire [63:0] T_6662;
  wire [63:0] GEN_700;
  wire [63:0] T_6663;
  wire [63:0] GEN_701;
  wire [63:0] T_6664;
  wire [63:0] T_6665;
  wire [63:0] T_6666;
  wire [63:0] T_6667;
  wire [63:0] T_6668;
  wire [63:0] T_6669;
  wire [63:0] T_6670;
  wire [63:0] T_6671;
  wire [63:0] GEN_702;
  wire [63:0] T_6672;
  wire [63:0] T_6673;
  wire [63:0] T_6674;
  wire [63:0] T_6675;
  wire [63:0] T_6676;
  wire [63:0] T_6677;
  wire [63:0] T_6678;
  wire [63:0] T_6679;
  wire [4:0] T_6680;
  wire [4:0] GEN_139;
  wire [1:0] supportedModes_0;
  wire [1:0] supportedModes_1;
  wire [1:0] supportedModes_2;
  wire  T_6738_debug;
  wire [1:0] T_6738_prv;
  wire  T_6738_sd;
  wire [30:0] T_6738_zero3;
  wire  T_6738_sd_rv32;
  wire [1:0] T_6738_zero2;
  wire [4:0] T_6738_vm;
  wire [4:0] T_6738_zero1;
  wire  T_6738_pum;
  wire  T_6738_mprv;
  wire [1:0] T_6738_xs;
  wire [1:0] T_6738_fs;
  wire [1:0] T_6738_mpp;
  wire [1:0] T_6738_hpp;
  wire  T_6738_spp;
  wire  T_6738_mpie;
  wire  T_6738_hpie;
  wire  T_6738_spie;
  wire  T_6738_upie;
  wire  T_6738_mie;
  wire  T_6738_hie;
  wire  T_6738_sie;
  wire  T_6738_uie;
  wire [66:0] T_6763;
  wire  T_6764;
  wire  T_6765;
  wire  T_6766;
  wire  T_6767;
  wire  T_6768;
  wire  T_6769;
  wire  T_6770;
  wire  T_6771;
  wire  T_6772;
  wire [1:0] T_6773;
  wire [1:0] T_6774;
  wire [1:0] T_6775;
  wire [1:0] T_6776;
  wire  T_6777;
  wire  T_6778;
  wire [4:0] T_6779;
  wire [4:0] T_6780;
  wire [1:0] T_6781;
  wire  T_6782;
  wire [30:0] T_6783;
  wire  T_6784;
  wire [1:0] T_6785;
  wire  T_6786;
  wire  T_6787;
  wire  T_6788;
  wire  T_6789;
  wire  T_6792;
  wire  T_6793;
  wire [1:0] GEN_140;
  wire [4:0] GEN_707;
  wire  T_6795;
  wire [4:0] GEN_141;
  wire [4:0] GEN_708;
  wire  T_6798;
  wire [4:0] GEN_142;
  wire  T_6801;
  wire [1:0] GEN_710;
  wire [2:0] T_6803;
  wire [1:0] T_6804;
  wire  GEN_167;
  wire  GEN_168;
  wire  GEN_169;
  wire [1:0] GEN_170;
  wire  GEN_171;
  wire [1:0] GEN_172;
  wire  GEN_173;
  wire  GEN_174;
  wire [4:0] GEN_175;
  wire [1:0] GEN_176;
  wire  T_6833_rocc;
  wire  T_6833_meip;
  wire  T_6833_heip;
  wire  T_6833_seip;
  wire  T_6833_ueip;
  wire  T_6833_mtip;
  wire  T_6833_htip;
  wire  T_6833_stip;
  wire  T_6833_utip;
  wire  T_6833_msip;
  wire  T_6833_hsip;
  wire  T_6833_ssip;
  wire  T_6833_usip;
  wire  T_6847;
  wire  T_6848;
  wire  T_6849;
  wire  T_6850;
  wire  T_6851;
  wire  T_6852;
  wire  T_6853;
  wire  T_6854;
  wire  T_6855;
  wire  T_6856;
  wire  T_6857;
  wire  T_6858;
  wire  T_6859;
  wire  GEN_190;
  wire  GEN_191;
  wire [63:0] GEN_711;
  wire [63:0] T_6860;
  wire [63:0] GEN_192;
  wire [63:0] T_6861;
  wire [63:0] T_6863;
  wire [63:0] T_6864;
  wire [63:0] GEN_193;
  wire [63:0] GEN_194;
  wire [61:0] T_6865;
  wire [63:0] GEN_713;
  wire [63:0] T_6866;
  wire [63:0] GEN_195;
  wire [63:0] T_6868;
  wire [63:0] GEN_196;
  wire [39:0] T_6869;
  wire [39:0] GEN_197;
  wire [1:0] T_6906_xdebugver;
  wire  T_6906_ndreset;
  wire  T_6906_fullreset;
  wire [11:0] T_6906_hwbpcount;
  wire  T_6906_ebreakm;
  wire  T_6906_ebreakh;
  wire  T_6906_ebreaks;
  wire  T_6906_ebreaku;
  wire  T_6906_zero2;
  wire  T_6906_stopcycle;
  wire  T_6906_stoptime;
  wire [2:0] T_6906_cause;
  wire  T_6906_debugint;
  wire  T_6906_zero1;
  wire  T_6906_halt;
  wire  T_6906_step;
  wire [1:0] T_6906_prv;
  wire [1:0] T_6924;
  wire [2:0] T_6929;
  wire  T_6934;
  wire  T_6935;
  wire  T_6936;
  wire [11:0] T_6937;
  wire  T_6938;
  wire  T_6939;
  wire [1:0] T_6940;
  wire  GEN_215;
  wire  GEN_216;
  wire  GEN_217;
  wire  GEN_218;
  wire  GEN_219;
  wire [1:0] GEN_220;
  wire [63:0] GEN_221;
  wire [63:0] GEN_222;
  wire  T_6993_debug;
  wire [1:0] T_6993_prv;
  wire  T_6993_sd;
  wire [30:0] T_6993_zero3;
  wire  T_6993_sd_rv32;
  wire [1:0] T_6993_zero2;
  wire [4:0] T_6993_vm;
  wire [4:0] T_6993_zero1;
  wire  T_6993_pum;
  wire  T_6993_mprv;
  wire [1:0] T_6993_xs;
  wire [1:0] T_6993_fs;
  wire [1:0] T_6993_mpp;
  wire [1:0] T_6993_hpp;
  wire  T_6993_spp;
  wire  T_6993_mpie;
  wire  T_6993_hpie;
  wire  T_6993_spie;
  wire  T_6993_upie;
  wire  T_6993_mie;
  wire  T_6993_hie;
  wire  T_6993_sie;
  wire  T_6993_uie;
  wire [66:0] T_7018;
  wire  T_7019;
  wire  T_7020;
  wire  T_7021;
  wire  T_7022;
  wire  T_7023;
  wire  T_7024;
  wire  T_7025;
  wire  T_7026;
  wire  T_7027;
  wire [1:0] T_7028;
  wire [1:0] T_7029;
  wire [1:0] T_7030;
  wire [1:0] T_7031;
  wire  T_7032;
  wire  T_7033;
  wire [4:0] T_7034;
  wire [4:0] T_7035;
  wire [1:0] T_7036;
  wire  T_7037;
  wire [30:0] T_7038;
  wire  T_7039;
  wire [1:0] T_7040;
  wire  T_7041;
  wire  T_7043;
  wire [1:0] GEN_716;
  wire [2:0] T_7045;
  wire [1:0] T_7046;
  wire  GEN_247;
  wire  GEN_248;
  wire [1:0] GEN_249;
  wire  GEN_250;
  wire [1:0] GEN_251;
  wire  T_7075_rocc;
  wire  T_7075_meip;
  wire  T_7075_heip;
  wire  T_7075_seip;
  wire  T_7075_ueip;
  wire  T_7075_mtip;
  wire  T_7075_htip;
  wire  T_7075_stip;
  wire  T_7075_utip;
  wire  T_7075_msip;
  wire  T_7075_hsip;
  wire  T_7075_ssip;
  wire  T_7075_usip;
  wire  GEN_265;
  wire [63:0] T_7103;
  wire [63:0] T_7104;
  wire [63:0] T_7105;
  wire [63:0] GEN_266;
  wire [63:0] GEN_267;
  wire [19:0] T_7106;
  wire [37:0] GEN_268;
  wire [63:0] GEN_269;
  wire [63:0] GEN_270;
  wire [63:0] GEN_271;
  wire [39:0] GEN_272;
  wire [63:0] GEN_719;
  wire [63:0] T_7114;
  wire [63:0] GEN_273;
  wire [63:0] GEN_720;
  wire [63:0] T_7115;
  wire [63:0] GEN_274;
  wire  T_7124_tdrmode;
  wire [61:0] T_7124_reserved;
  wire  T_7124_tdrindex;
  wire [61:0] T_7129;
  wire  T_7130;
  wire  GEN_275;
  wire  T_7131;
  wire [3:0] T_7158_tdrtype;
  wire [4:0] T_7158_bpamaskmax;
  wire [35:0] T_7158_reserved;
  wire [7:0] T_7158_bpaction;
  wire [3:0] T_7158_bpmatch;
  wire  T_7158_m;
  wire  T_7158_h;
  wire  T_7158_s;
  wire  T_7158_u;
  wire  T_7158_r;
  wire  T_7158_w;
  wire  T_7158_x;
  wire [3:0] T_7178;
  wire [7:0] T_7179;
  wire [35:0] T_7180;
  wire [4:0] T_7181;
  wire [3:0] T_7182;
  wire [3:0] GEN_13;
  wire [4:0] GEN_14;
  wire [35:0] GEN_15;
  wire [7:0] GEN_16;
  wire [3:0] GEN_17;
  wire [3:0] GEN_284;
  wire  GEN_18;
  wire  GEN_286;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_290;
  wire  GEN_21;
  wire  GEN_292;
  wire  GEN_22;
  wire  GEN_294;
  wire  GEN_23;
  wire  GEN_296;
  wire  GEN_24;
  wire  GEN_298;
  wire [3:0] GEN_721;
  wire [3:0] T_7212;
  wire [3:0] GEN_25;
  wire [3:0] GEN_300;
  wire [3:0] GEN_327;
  wire  GEN_330;
  wire  GEN_336;
  wire  GEN_339;
  wire  GEN_342;
  wire  GEN_345;
  wire  GEN_348;
  wire [38:0] GEN_26;
  wire [38:0] GEN_351;
  wire [38:0] GEN_354;
  wire [3:0] GEN_381;
  wire  GEN_384;
  wire  GEN_390;
  wire  GEN_393;
  wire  GEN_396;
  wire  GEN_399;
  wire  GEN_402;
  wire [38:0] GEN_406;
  wire  GEN_432;
  wire  GEN_433;
  wire  GEN_434;
  wire [1:0] GEN_435;
  wire  GEN_436;
  wire [1:0] GEN_437;
  wire  GEN_438;
  wire  GEN_439;
  wire [4:0] GEN_440;
  wire [1:0] GEN_441;
  wire  GEN_455;
  wire  GEN_456;
  wire [63:0] GEN_457;
  wire [63:0] GEN_458;
  wire [63:0] GEN_459;
  wire [63:0] GEN_460;
  wire [63:0] GEN_461;
  wire [39:0] GEN_462;
  wire  GEN_480;
  wire  GEN_481;
  wire  GEN_482;
  wire  GEN_483;
  wire  GEN_484;
  wire [1:0] GEN_485;
  wire [63:0] GEN_486;
  wire [63:0] GEN_487;
  wire [63:0] GEN_525;
  wire [37:0] GEN_526;
  wire [63:0] GEN_527;
  wire [63:0] GEN_528;
  wire [63:0] GEN_529;
  wire [39:0] GEN_530;
  wire [63:0] GEN_531;
  wire [63:0] GEN_532;
  wire  GEN_536;
  wire [3:0] GEN_562;
  wire  GEN_565;
  wire  GEN_571;
  wire  GEN_574;
  wire  GEN_577;
  wire  GEN_580;
  wire  GEN_583;
  wire [38:0] GEN_587;
  wire  GEN_589;
  wire  GEN_590;
  wire  GEN_591;
  wire [3:0] T_7278_control_tdrtype;
  wire [4:0] T_7278_control_bpamaskmax;
  wire [35:0] T_7278_control_reserved;
  wire [7:0] T_7278_control_bpaction;
  wire [3:0] T_7278_control_bpmatch;
  wire  T_7278_control_m;
  wire  T_7278_control_h;
  wire  T_7278_control_s;
  wire  T_7278_control_u;
  wire  T_7278_control_r;
  wire  T_7278_control_w;
  wire  T_7278_control_x;
  wire [38:0] T_7278_address;
  wire [102:0] T_7294;
  wire [38:0] T_7295;
  wire  T_7296;
  wire  T_7297;
  wire  T_7298;
  wire  T_7299;
  wire  T_7300;
  wire  T_7301;
  wire  T_7302;
  wire [3:0] T_7303;
  wire [7:0] T_7304;
  wire [35:0] T_7305;
  wire [4:0] T_7306;
  wire [3:0] T_7307;
  reg  GEN_63;
  reg [31:0] GEN_416;
  reg [6:0] GEN_143;
  reg [31:0] GEN_417;
  reg [4:0] GEN_144;
  reg [31:0] GEN_418;
  reg [4:0] GEN_145;
  reg [31:0] GEN_419;
  reg  GEN_146;
  reg [31:0] GEN_420;
  reg  GEN_147;
  reg [31:0] GEN_421;
  reg  GEN_148;
  reg [31:0] GEN_422;
  reg [4:0] GEN_149;
  reg [31:0] GEN_423;
  reg [6:0] GEN_150;
  reg [31:0] GEN_424;
  reg [63:0] GEN_151;
  reg [63:0] GEN_425;
  reg [63:0] GEN_152;
  reg [63:0] GEN_426;
  reg  GEN_153;
  reg [31:0] GEN_427;
  reg  GEN_154;
  reg [31:0] GEN_428;
  reg  GEN_155;
  reg [31:0] GEN_429;
  reg  GEN_156;
  reg [31:0] GEN_430;
  reg [39:0] GEN_157;
  reg [63:0] GEN_431;
  reg [8:0] GEN_158;
  reg [31:0] GEN_442;
  reg [4:0] GEN_159;
  reg [31:0] GEN_443;
  reg [2:0] GEN_160;
  reg [31:0] GEN_444;
  reg [63:0] GEN_161;
  reg [63:0] GEN_445;
  reg  GEN_162;
  reg [31:0] GEN_446;
  reg  GEN_163;
  reg [31:0] GEN_447;
  reg [63:0] GEN_164;
  reg [63:0] GEN_448;
  reg [63:0] GEN_165;
  reg [63:0] GEN_449;
  reg  GEN_166;
  reg [31:0] GEN_450;
  reg  GEN_177;
  reg [31:0] GEN_451;
  reg  GEN_178;
  reg [31:0] GEN_452;
  reg  GEN_179;
  reg [31:0] GEN_453;
  reg  GEN_180;
  reg [31:0] GEN_454;
  reg  GEN_181;
  reg [31:0] GEN_463;
  reg  GEN_182;
  reg [31:0] GEN_464;
  reg [1:0] GEN_183;
  reg [31:0] GEN_465;
  reg  GEN_184;
  reg [31:0] GEN_466;
  reg [30:0] GEN_185;
  reg [31:0] GEN_467;
  reg  GEN_186;
  reg [31:0] GEN_468;
  reg [1:0] GEN_187;
  reg [31:0] GEN_469;
  reg [4:0] GEN_188;
  reg [31:0] GEN_470;
  reg [4:0] GEN_189;
  reg [31:0] GEN_471;
  reg  GEN_198;
  reg [31:0] GEN_472;
  reg  GEN_199;
  reg [31:0] GEN_473;
  reg [1:0] GEN_200;
  reg [31:0] GEN_474;
  reg [1:0] GEN_201;
  reg [31:0] GEN_475;
  reg [1:0] GEN_202;
  reg [31:0] GEN_476;
  reg [1:0] GEN_203;
  reg [31:0] GEN_477;
  reg  GEN_204;
  reg [31:0] GEN_478;
  reg  GEN_205;
  reg [31:0] GEN_479;
  reg  GEN_206;
  reg [31:0] GEN_488;
  reg  GEN_207;
  reg [31:0] GEN_489;
  reg  GEN_208;
  reg [31:0] GEN_490;
  reg  GEN_209;
  reg [31:0] GEN_491;
  reg  GEN_210;
  reg [31:0] GEN_492;
  reg  GEN_211;
  reg [31:0] GEN_493;
  reg  GEN_212;
  reg [31:0] GEN_494;
  reg  GEN_213;
  reg [31:0] GEN_495;
  reg  GEN_214;
  reg [31:0] GEN_496;
  reg [2:0] GEN_223;
  reg [31:0] GEN_497;
  reg [1:0] GEN_224;
  reg [31:0] GEN_498;
  reg [2:0] GEN_225;
  reg [31:0] GEN_499;
  reg  GEN_226;
  reg [31:0] GEN_500;
  reg [3:0] GEN_227;
  reg [31:0] GEN_501;
  reg [63:0] GEN_228;
  reg [63:0] GEN_502;
  reg  GEN_229;
  reg [31:0] GEN_503;
  reg  GEN_230;
  reg [31:0] GEN_504;
  reg [64:0] GEN_231;
  reg [95:0] GEN_505;
  reg [4:0] GEN_232;
  reg [31:0] GEN_506;
  reg  GEN_233;
  reg [31:0] GEN_507;
  reg  GEN_234;
  reg [31:0] GEN_508;
  assign io_rw_rdata = T_6679;
  assign io_csr_stall = reg_wfi;
  assign io_csr_xcpt = T_6436;
  assign io_eret = insn_ret;
  assign io_singleStep = T_6488;
  assign io_status_debug = reg_debug;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_sd = T_6495;
  assign io_status_zero3 = reg_mstatus_zero3;
  assign io_status_sd_rv32 = reg_mstatus_sd_rv32;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign io_status_vm = reg_mstatus_vm;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign io_status_pum = reg_mstatus_pum;
  assign io_status_mprv = reg_mstatus_mprv;
  assign io_status_xs = reg_mstatus_xs;
  assign io_status_fs = reg_mstatus_fs;
  assign io_status_mpp = reg_mstatus_mpp;
  assign io_status_hpp = reg_mstatus_hpp;
  assign io_status_spp = reg_mstatus_spp;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_hpie = reg_mstatus_hpie;
  assign io_status_spie = reg_mstatus_spie;
  assign io_status_upie = reg_mstatus_upie;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = reg_mstatus_hie;
  assign io_status_sie = reg_mstatus_sie;
  assign io_status_uie = reg_mstatus_uie;
  assign io_ptbr_asid = reg_sptbr_asid;
  assign io_ptbr_ppn = reg_sptbr_ppn;
  assign io_evec = T_6485;
  assign io_fatc = insn_sfence_vm;
  assign io_time = reg_cycle;
  assign io_fcsr_rm = reg_frm;
  assign io_rocc_cmd_valid = GEN_63;
  assign io_rocc_cmd_bits_inst_funct = GEN_143;
  assign io_rocc_cmd_bits_inst_rs2 = GEN_144;
  assign io_rocc_cmd_bits_inst_rs1 = GEN_145;
  assign io_rocc_cmd_bits_inst_xd = GEN_146;
  assign io_rocc_cmd_bits_inst_xs1 = GEN_147;
  assign io_rocc_cmd_bits_inst_xs2 = GEN_148;
  assign io_rocc_cmd_bits_inst_rd = GEN_149;
  assign io_rocc_cmd_bits_inst_opcode = GEN_150;
  assign io_rocc_cmd_bits_rs1 = GEN_151;
  assign io_rocc_cmd_bits_rs2 = GEN_152;
  assign io_rocc_resp_ready = GEN_153;
  assign io_rocc_mem_req_ready = GEN_154;
  assign io_rocc_mem_s2_nack = GEN_155;
  assign io_rocc_mem_resp_valid = GEN_156;
  assign io_rocc_mem_resp_bits_addr = GEN_157;
  assign io_rocc_mem_resp_bits_tag = GEN_158;
  assign io_rocc_mem_resp_bits_cmd = GEN_159;
  assign io_rocc_mem_resp_bits_typ = GEN_160;
  assign io_rocc_mem_resp_bits_data = GEN_161;
  assign io_rocc_mem_resp_bits_replay = GEN_162;
  assign io_rocc_mem_resp_bits_has_data = GEN_163;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_164;
  assign io_rocc_mem_resp_bits_store_data = GEN_165;
  assign io_rocc_mem_replay_next = GEN_166;
  assign io_rocc_mem_xcpt_ma_ld = GEN_177;
  assign io_rocc_mem_xcpt_ma_st = GEN_178;
  assign io_rocc_mem_xcpt_pf_ld = GEN_179;
  assign io_rocc_mem_xcpt_pf_st = GEN_180;
  assign io_rocc_mem_ordered = GEN_181;
  assign io_rocc_status_debug = GEN_182;
  assign io_rocc_status_prv = GEN_183;
  assign io_rocc_status_sd = GEN_184;
  assign io_rocc_status_zero3 = GEN_185;
  assign io_rocc_status_sd_rv32 = GEN_186;
  assign io_rocc_status_zero2 = GEN_187;
  assign io_rocc_status_vm = GEN_188;
  assign io_rocc_status_zero1 = GEN_189;
  assign io_rocc_status_pum = GEN_198;
  assign io_rocc_status_mprv = GEN_199;
  assign io_rocc_status_xs = GEN_200;
  assign io_rocc_status_fs = GEN_201;
  assign io_rocc_status_mpp = GEN_202;
  assign io_rocc_status_hpp = GEN_203;
  assign io_rocc_status_spp = GEN_204;
  assign io_rocc_status_mpie = GEN_205;
  assign io_rocc_status_hpie = GEN_206;
  assign io_rocc_status_spie = GEN_207;
  assign io_rocc_status_upie = GEN_208;
  assign io_rocc_status_mie = GEN_209;
  assign io_rocc_status_hie = GEN_210;
  assign io_rocc_status_sie = GEN_211;
  assign io_rocc_status_uie = GEN_212;
  assign io_rocc_autl_acquire_ready = GEN_213;
  assign io_rocc_autl_grant_valid = GEN_214;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_223;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_224;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_225;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_226;
  assign io_rocc_autl_grant_bits_g_type = GEN_227;
  assign io_rocc_autl_grant_bits_data = GEN_228;
  assign io_rocc_fpu_req_ready = GEN_229;
  assign io_rocc_fpu_resp_valid = GEN_230;
  assign io_rocc_fpu_resp_bits_data = GEN_231;
  assign io_rocc_fpu_resp_bits_exc = GEN_232;
  assign io_rocc_exception = GEN_233;
  assign io_rocc_csr_waddr = io_rw_addr;
  assign io_rocc_csr_wdata = wdata;
  assign io_rocc_csr_wen = wen;
  assign io_rocc_host_id = GEN_234;
  assign io_interrupt = GEN_65;
  assign io_interrupt_cause = GEN_66;
  assign io_bp_0_control_tdrtype = reg_bp_0_control_tdrtype;
  assign io_bp_0_control_bpamaskmax = reg_bp_0_control_bpamaskmax;
  assign io_bp_0_control_reserved = reg_bp_0_control_reserved;
  assign io_bp_0_control_bpaction = reg_bp_0_control_bpaction;
  assign io_bp_0_control_bpmatch = reg_bp_0_control_bpmatch;
  assign io_bp_0_control_m = reg_bp_0_control_m;
  assign io_bp_0_control_h = reg_bp_0_control_h;
  assign io_bp_0_control_s = reg_bp_0_control_s;
  assign io_bp_0_control_u = reg_bp_0_control_u;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_bp_0_address = reg_bp_0_address;
  assign T_4992_debug = T_5040;
  assign T_4992_prv = T_5039;
  assign T_4992_sd = T_5038;
  assign T_4992_zero3 = T_5037;
  assign T_4992_sd_rv32 = T_5036;
  assign T_4992_zero2 = T_5035;
  assign T_4992_vm = T_5034;
  assign T_4992_zero1 = T_5033;
  assign T_4992_pum = T_5032;
  assign T_4992_mprv = T_5031;
  assign T_4992_xs = T_5030;
  assign T_4992_fs = T_5029;
  assign T_4992_mpp = T_5028;
  assign T_4992_hpp = T_5027;
  assign T_4992_spp = T_5026;
  assign T_4992_mpie = T_5025;
  assign T_4992_hpie = T_5024;
  assign T_4992_spie = T_5023;
  assign T_4992_upie = T_5022;
  assign T_4992_mie = T_5021;
  assign T_4992_hie = T_5020;
  assign T_4992_sie = T_5019;
  assign T_4992_uie = T_5018;
  assign T_5017 = {{66'd0}, 1'h0};
  assign T_5018 = T_5017[0];
  assign T_5019 = T_5017[1];
  assign T_5020 = T_5017[2];
  assign T_5021 = T_5017[3];
  assign T_5022 = T_5017[4];
  assign T_5023 = T_5017[5];
  assign T_5024 = T_5017[6];
  assign T_5025 = T_5017[7];
  assign T_5026 = T_5017[8];
  assign T_5027 = T_5017[10:9];
  assign T_5028 = T_5017[12:11];
  assign T_5029 = T_5017[14:13];
  assign T_5030 = T_5017[16:15];
  assign T_5031 = T_5017[17];
  assign T_5032 = T_5017[18];
  assign T_5033 = T_5017[23:19];
  assign T_5034 = T_5017[28:24];
  assign T_5035 = T_5017[30:29];
  assign T_5036 = T_5017[31];
  assign T_5037 = T_5017[62:32];
  assign T_5038 = T_5017[63];
  assign T_5039 = T_5017[65:64];
  assign T_5040 = T_5017[66];
  assign reset_mstatus_debug = T_4992_debug;
  assign reset_mstatus_prv = 2'h3;
  assign reset_mstatus_sd = T_4992_sd;
  assign reset_mstatus_zero3 = T_4992_zero3;
  assign reset_mstatus_sd_rv32 = T_4992_sd_rv32;
  assign reset_mstatus_zero2 = T_4992_zero2;
  assign reset_mstatus_vm = T_4992_vm;
  assign reset_mstatus_zero1 = T_4992_zero1;
  assign reset_mstatus_pum = T_4992_pum;
  assign reset_mstatus_mprv = T_4992_mprv;
  assign reset_mstatus_xs = T_4992_xs;
  assign reset_mstatus_fs = T_4992_fs;
  assign reset_mstatus_mpp = 2'h3;
  assign reset_mstatus_hpp = T_4992_hpp;
  assign reset_mstatus_spp = T_4992_spp;
  assign reset_mstatus_mpie = T_4992_mpie;
  assign reset_mstatus_hpie = T_4992_hpie;
  assign reset_mstatus_spie = T_4992_spie;
  assign reset_mstatus_upie = T_4992_upie;
  assign reset_mstatus_mie = T_4992_mie;
  assign reset_mstatus_hie = T_4992_hie;
  assign reset_mstatus_sie = T_4992_sie;
  assign reset_mstatus_uie = T_4992_uie;
  assign T_5126_xdebugver = T_5162;
  assign T_5126_ndreset = T_5161;
  assign T_5126_fullreset = T_5160;
  assign T_5126_hwbpcount = T_5159;
  assign T_5126_ebreakm = T_5158;
  assign T_5126_ebreakh = T_5157;
  assign T_5126_ebreaks = T_5156;
  assign T_5126_ebreaku = T_5155;
  assign T_5126_zero2 = T_5154;
  assign T_5126_stopcycle = T_5153;
  assign T_5126_stoptime = T_5152;
  assign T_5126_cause = T_5151;
  assign T_5126_debugint = T_5150;
  assign T_5126_zero1 = T_5149;
  assign T_5126_halt = T_5148;
  assign T_5126_step = T_5147;
  assign T_5126_prv = T_5146;
  assign T_5145 = {{31'd0}, 1'h0};
  assign T_5146 = T_5145[1:0];
  assign T_5147 = T_5145[2];
  assign T_5148 = T_5145[3];
  assign T_5149 = T_5145[4];
  assign T_5150 = T_5145[5];
  assign T_5151 = T_5145[8:6];
  assign T_5152 = T_5145[9];
  assign T_5153 = T_5145[10];
  assign T_5154 = T_5145[11];
  assign T_5155 = T_5145[12];
  assign T_5156 = T_5145[13];
  assign T_5157 = T_5145[14];
  assign T_5158 = T_5145[15];
  assign T_5159 = T_5145[27:16];
  assign T_5160 = T_5145[28];
  assign T_5161 = T_5145[29];
  assign T_5162 = T_5145[31:30];
  assign reset_dcsr_xdebugver = {{1'd0}, 1'h1};
  assign reset_dcsr_ndreset = T_5126_ndreset;
  assign reset_dcsr_fullreset = T_5126_fullreset;
  assign reset_dcsr_hwbpcount = T_5126_hwbpcount;
  assign reset_dcsr_ebreakm = T_5126_ebreakm;
  assign reset_dcsr_ebreakh = T_5126_ebreakh;
  assign reset_dcsr_ebreaks = T_5126_ebreaks;
  assign reset_dcsr_ebreaku = T_5126_ebreaku;
  assign reset_dcsr_zero2 = T_5126_zero2;
  assign reset_dcsr_stopcycle = T_5126_stopcycle;
  assign reset_dcsr_stoptime = T_5126_stoptime;
  assign reset_dcsr_cause = T_5126_cause;
  assign reset_dcsr_debugint = T_5126_debugint;
  assign reset_dcsr_zero1 = T_5126_zero1;
  assign reset_dcsr_halt = T_5126_halt;
  assign reset_dcsr_step = T_5126_step;
  assign reset_dcsr_prv = 2'h3;
  assign T_5228_rocc = T_5256;
  assign T_5228_meip = T_5255;
  assign T_5228_heip = T_5254;
  assign T_5228_seip = T_5253;
  assign T_5228_ueip = T_5252;
  assign T_5228_mtip = T_5251;
  assign T_5228_htip = T_5250;
  assign T_5228_stip = T_5249;
  assign T_5228_utip = T_5248;
  assign T_5228_msip = T_5247;
  assign T_5228_hsip = T_5246;
  assign T_5228_ssip = T_5245;
  assign T_5228_usip = T_5244;
  assign T_5243 = {{12'd0}, 1'h0};
  assign T_5244 = T_5243[0];
  assign T_5245 = T_5243[1];
  assign T_5246 = T_5243[2];
  assign T_5247 = T_5243[3];
  assign T_5248 = T_5243[4];
  assign T_5249 = T_5243[5];
  assign T_5250 = T_5243[6];
  assign T_5251 = T_5243[7];
  assign T_5252 = T_5243[8];
  assign T_5253 = T_5243[9];
  assign T_5254 = T_5243[10];
  assign T_5255 = T_5243[11];
  assign T_5256 = T_5243[12];
  assign T_5257_rocc = 1'h0;
  assign T_5257_meip = 1'h1;
  assign T_5257_heip = T_5228_heip;
  assign T_5257_seip = 1'h1;
  assign T_5257_ueip = T_5228_ueip;
  assign T_5257_mtip = 1'h1;
  assign T_5257_htip = T_5228_htip;
  assign T_5257_stip = 1'h1;
  assign T_5257_utip = T_5228_utip;
  assign T_5257_msip = 1'h1;
  assign T_5257_hsip = T_5228_hsip;
  assign T_5257_ssip = 1'h1;
  assign T_5257_usip = T_5228_usip;
  assign T_5278_rocc = T_5257_rocc;
  assign T_5278_meip = 1'h0;
  assign T_5278_heip = T_5257_heip;
  assign T_5278_seip = T_5257_seip;
  assign T_5278_ueip = T_5257_ueip;
  assign T_5278_mtip = 1'h0;
  assign T_5278_htip = T_5257_htip;
  assign T_5278_stip = T_5257_stip;
  assign T_5278_utip = T_5257_utip;
  assign T_5278_msip = 1'h0;
  assign T_5278_hsip = T_5257_hsip;
  assign T_5278_ssip = T_5257_ssip;
  assign T_5278_usip = T_5257_usip;
  assign T_5295 = {T_5257_hsip,T_5257_ssip};
  assign T_5296 = {T_5295,T_5257_usip};
  assign T_5297 = {T_5257_stip,T_5257_utip};
  assign T_5298 = {T_5297,T_5257_msip};
  assign T_5299 = {T_5298,T_5296};
  assign T_5300 = {T_5257_ueip,T_5257_mtip};
  assign T_5301 = {T_5300,T_5257_htip};
  assign T_5302 = {T_5257_heip,T_5257_seip};
  assign T_5303 = {T_5257_rocc,T_5257_meip};
  assign T_5304 = {T_5303,T_5302};
  assign T_5305 = {T_5304,T_5301};
  assign supported_interrupts = {T_5305,T_5299};
  assign T_5306 = {T_5278_hsip,T_5278_ssip};
  assign T_5307 = {T_5306,T_5278_usip};
  assign T_5308 = {T_5278_stip,T_5278_utip};
  assign T_5309 = {T_5308,T_5278_msip};
  assign T_5310 = {T_5309,T_5307};
  assign T_5311 = {T_5278_ueip,T_5278_mtip};
  assign T_5312 = {T_5311,T_5278_htip};
  assign T_5313 = {T_5278_heip,T_5278_seip};
  assign T_5314 = {T_5278_rocc,T_5278_meip};
  assign T_5315 = {T_5314,T_5313};
  assign T_5316 = {T_5315,T_5312};
  assign delegable_interrupts = {T_5316,T_5310};
  assign exception = io_exception | io_csr_xcpt;
  assign T_5322 = io_retire | exception;
  assign GEN_27 = T_5322 ? 1'h1 : reg_singleStepped;
  assign T_5325 = io_singleStep == 1'h0;
  assign GEN_28 = T_5325 ? 1'h0 : GEN_27;
  assign T_5336 = reg_singleStepped == 1'h0;
  assign T_5338 = io_retire == 1'h0;
  assign T_5339 = T_5336 | T_5338;
  assign T_5340 = T_5339 | reset;
  assign T_5342 = T_5340 == 1'h0;
  assign GEN_595 = {{1'd0}, T_5544};
  assign T_5548 = GEN_595 + 7'h1;
  assign T_5549 = T_5548[6:0];
  assign T_5550 = T_5549[5:0];
  assign GEN_29 = io_uarch_counters_0 ? T_5550 : T_5544;
  assign T_5553 = T_5549[6];
  assign T_5554 = io_uarch_counters_0 & T_5553;
  assign GEN_596 = {{57'd0}, 1'h1};
  assign T_5556 = T_5552 + GEN_596;
  assign T_5557 = T_5556[57:0];
  assign GEN_30 = T_5554 ? T_5557 : T_5552;
  assign GEN_597 = {{1'd0}, T_5560};
  assign T_5564 = GEN_597 + 7'h1;
  assign T_5565 = T_5564[6:0];
  assign T_5566 = T_5565[5:0];
  assign GEN_31 = io_uarch_counters_1 ? T_5566 : T_5560;
  assign T_5569 = T_5565[6];
  assign T_5570 = io_uarch_counters_1 & T_5569;
  assign T_5572 = T_5568 + GEN_596;
  assign T_5573 = T_5572[57:0];
  assign GEN_32 = T_5570 ? T_5573 : T_5568;
  assign GEN_599 = {{1'd0}, T_5576};
  assign T_5580 = GEN_599 + 7'h1;
  assign T_5581 = T_5580[6:0];
  assign T_5582 = T_5581[5:0];
  assign GEN_33 = io_uarch_counters_2 ? T_5582 : T_5576;
  assign T_5585 = T_5581[6];
  assign T_5586 = io_uarch_counters_2 & T_5585;
  assign T_5588 = T_5584 + GEN_596;
  assign T_5589 = T_5588[57:0];
  assign GEN_34 = T_5586 ? T_5589 : T_5584;
  assign GEN_601 = {{1'd0}, T_5592};
  assign T_5596 = GEN_601 + 7'h1;
  assign T_5597 = T_5596[6:0];
  assign T_5598 = T_5597[5:0];
  assign GEN_35 = io_uarch_counters_3 ? T_5598 : T_5592;
  assign T_5601 = T_5597[6];
  assign T_5602 = io_uarch_counters_3 & T_5601;
  assign T_5604 = T_5600 + GEN_596;
  assign T_5605 = T_5604[57:0];
  assign GEN_36 = T_5602 ? T_5605 : T_5600;
  assign GEN_603 = {{1'd0}, T_5608};
  assign T_5612 = GEN_603 + 7'h1;
  assign T_5613 = T_5612[6:0];
  assign T_5614 = T_5613[5:0];
  assign GEN_37 = io_uarch_counters_4 ? T_5614 : T_5608;
  assign T_5617 = T_5613[6];
  assign T_5618 = io_uarch_counters_4 & T_5617;
  assign T_5620 = T_5616 + GEN_596;
  assign T_5621 = T_5620[57:0];
  assign GEN_38 = T_5618 ? T_5621 : T_5616;
  assign GEN_605 = {{1'd0}, T_5624};
  assign T_5628 = GEN_605 + 7'h1;
  assign T_5629 = T_5628[6:0];
  assign T_5630 = T_5629[5:0];
  assign GEN_39 = io_uarch_counters_5 ? T_5630 : T_5624;
  assign T_5633 = T_5629[6];
  assign T_5634 = io_uarch_counters_5 & T_5633;
  assign T_5636 = T_5632 + GEN_596;
  assign T_5637 = T_5636[57:0];
  assign GEN_40 = T_5634 ? T_5637 : T_5632;
  assign GEN_607 = {{1'd0}, T_5640};
  assign T_5644 = GEN_607 + 7'h1;
  assign T_5645 = T_5644[6:0];
  assign T_5646 = T_5645[5:0];
  assign GEN_41 = io_uarch_counters_6 ? T_5646 : T_5640;
  assign T_5649 = T_5645[6];
  assign T_5650 = io_uarch_counters_6 & T_5649;
  assign T_5652 = T_5648 + GEN_596;
  assign T_5653 = T_5652[57:0];
  assign GEN_42 = T_5650 ? T_5653 : T_5648;
  assign GEN_609 = {{1'd0}, T_5656};
  assign T_5660 = GEN_609 + 7'h1;
  assign T_5661 = T_5660[6:0];
  assign T_5662 = T_5661[5:0];
  assign GEN_43 = io_uarch_counters_7 ? T_5662 : T_5656;
  assign T_5665 = T_5661[6];
  assign T_5666 = io_uarch_counters_7 & T_5665;
  assign T_5668 = T_5664 + GEN_596;
  assign T_5669 = T_5668[57:0];
  assign GEN_44 = T_5666 ? T_5669 : T_5664;
  assign GEN_611 = {{1'd0}, T_5672};
  assign T_5676 = GEN_611 + 7'h1;
  assign T_5677 = T_5676[6:0];
  assign T_5678 = T_5677[5:0];
  assign GEN_45 = io_uarch_counters_8 ? T_5678 : T_5672;
  assign T_5681 = T_5677[6];
  assign T_5682 = io_uarch_counters_8 & T_5681;
  assign T_5684 = T_5680 + GEN_596;
  assign T_5685 = T_5684[57:0];
  assign GEN_46 = T_5682 ? T_5685 : T_5680;
  assign GEN_613 = {{1'd0}, T_5688};
  assign T_5692 = GEN_613 + 7'h1;
  assign T_5693 = T_5692[6:0];
  assign T_5694 = T_5693[5:0];
  assign GEN_47 = io_uarch_counters_9 ? T_5694 : T_5688;
  assign T_5697 = T_5693[6];
  assign T_5698 = io_uarch_counters_9 & T_5697;
  assign T_5700 = T_5696 + GEN_596;
  assign T_5701 = T_5700[57:0];
  assign GEN_48 = T_5698 ? T_5701 : T_5696;
  assign GEN_615 = {{1'd0}, T_5704};
  assign T_5708 = GEN_615 + 7'h1;
  assign T_5709 = T_5708[6:0];
  assign T_5710 = T_5709[5:0];
  assign GEN_49 = io_uarch_counters_10 ? T_5710 : T_5704;
  assign T_5713 = T_5709[6];
  assign T_5714 = io_uarch_counters_10 & T_5713;
  assign T_5716 = T_5712 + GEN_596;
  assign T_5717 = T_5716[57:0];
  assign GEN_50 = T_5714 ? T_5717 : T_5712;
  assign GEN_617 = {{1'd0}, T_5720};
  assign T_5724 = GEN_617 + 7'h1;
  assign T_5725 = T_5724[6:0];
  assign T_5726 = T_5725[5:0];
  assign GEN_51 = io_uarch_counters_11 ? T_5726 : T_5720;
  assign T_5729 = T_5725[6];
  assign T_5730 = io_uarch_counters_11 & T_5729;
  assign T_5732 = T_5728 + GEN_596;
  assign T_5733 = T_5732[57:0];
  assign GEN_52 = T_5730 ? T_5733 : T_5728;
  assign GEN_619 = {{1'd0}, T_5736};
  assign T_5740 = GEN_619 + 7'h1;
  assign T_5741 = T_5740[6:0];
  assign T_5742 = T_5741[5:0];
  assign GEN_53 = io_uarch_counters_12 ? T_5742 : T_5736;
  assign T_5745 = T_5741[6];
  assign T_5746 = io_uarch_counters_12 & T_5745;
  assign T_5748 = T_5744 + GEN_596;
  assign T_5749 = T_5748[57:0];
  assign GEN_54 = T_5746 ? T_5749 : T_5744;
  assign GEN_621 = {{1'd0}, T_5752};
  assign T_5756 = GEN_621 + 7'h1;
  assign T_5757 = T_5756[6:0];
  assign T_5758 = T_5757[5:0];
  assign GEN_55 = io_uarch_counters_13 ? T_5758 : T_5752;
  assign T_5761 = T_5757[6];
  assign T_5762 = io_uarch_counters_13 & T_5761;
  assign T_5764 = T_5760 + GEN_596;
  assign T_5765 = T_5764[57:0];
  assign GEN_56 = T_5762 ? T_5765 : T_5760;
  assign GEN_623 = {{1'd0}, T_5768};
  assign T_5772 = GEN_623 + 7'h1;
  assign T_5773 = T_5772[6:0];
  assign T_5774 = T_5773[5:0];
  assign GEN_57 = io_uarch_counters_14 ? T_5774 : T_5768;
  assign T_5777 = T_5773[6];
  assign T_5778 = io_uarch_counters_14 & T_5777;
  assign T_5780 = T_5776 + GEN_596;
  assign T_5781 = T_5780[57:0];
  assign GEN_58 = T_5778 ? T_5781 : T_5776;
  assign GEN_625 = {{1'd0}, T_5784};
  assign T_5788 = GEN_625 + 7'h1;
  assign T_5789 = T_5788[6:0];
  assign T_5790 = T_5789[5:0];
  assign GEN_59 = io_uarch_counters_15 ? T_5790 : T_5784;
  assign T_5793 = T_5789[6];
  assign T_5794 = io_uarch_counters_15 & T_5793;
  assign T_5796 = T_5792 + GEN_596;
  assign T_5797 = T_5796[57:0];
  assign GEN_60 = T_5794 ? T_5797 : T_5792;
  assign GEN_627 = {{1'd0}, T_5802};
  assign T_5806 = GEN_627 + 7'h1;
  assign T_5807 = T_5806[6:0];
  assign T_5808 = T_5807[5:0];
  assign GEN_61 = io_retire ? T_5808 : T_5802;
  assign T_5811 = T_5807[6];
  assign T_5812 = io_retire & T_5811;
  assign T_5814 = T_5810 + GEN_596;
  assign T_5815 = T_5814[57:0];
  assign GEN_62 = T_5812 ? T_5815 : T_5810;
  assign T_5816 = {T_5810,T_5802};
  assign GEN_629 = {{1'd0}, T_5819};
  assign T_5823 = GEN_629 + 7'h1;
  assign T_5824 = T_5823[6:0];
  assign T_5825 = T_5824[5:0];
  assign T_5828 = T_5824[6];
  assign T_5831 = T_5827 + GEN_596;
  assign T_5832 = T_5831[57:0];
  assign GEN_64 = T_5828 ? T_5832 : T_5827;
  assign reg_cycle = {T_5827,T_5819};
  assign mip_rocc = io_rocc_interrupt;
  assign mip_meip = reg_mip_meip;
  assign mip_heip = reg_mip_heip;
  assign mip_seip = reg_mip_seip;
  assign mip_ueip = reg_mip_ueip;
  assign mip_mtip = reg_mip_mtip;
  assign mip_htip = reg_mip_htip;
  assign mip_stip = reg_mip_stip;
  assign mip_utip = reg_mip_utip;
  assign mip_msip = reg_mip_msip;
  assign mip_hsip = reg_mip_hsip;
  assign mip_ssip = reg_mip_ssip;
  assign mip_usip = reg_mip_usip;
  assign T_5846 = {mip_hsip,mip_ssip};
  assign T_5847 = {T_5846,mip_usip};
  assign T_5848 = {mip_stip,mip_utip};
  assign T_5849 = {T_5848,mip_msip};
  assign T_5850 = {T_5849,T_5847};
  assign T_5851 = {mip_ueip,mip_mtip};
  assign T_5852 = {T_5851,mip_htip};
  assign T_5853 = {mip_heip,mip_seip};
  assign T_5854 = {mip_rocc,mip_meip};
  assign T_5855 = {T_5854,T_5853};
  assign T_5856 = {T_5855,T_5852};
  assign T_5857 = {T_5856,T_5850};
  assign read_mip = T_5857 & supported_interrupts;
  assign GEN_631 = {{51'd0}, read_mip};
  assign pending_interrupts = GEN_631 & reg_mie;
  assign T_5859 = reg_debug == 1'h0;
  assign T_5861 = reg_mstatus_prv < 2'h3;
  assign T_5863 = reg_mstatus_prv == 2'h3;
  assign T_5864 = T_5863 & reg_mstatus_mie;
  assign T_5865 = T_5861 | T_5864;
  assign T_5866 = T_5859 & T_5865;
  assign T_5867 = ~ reg_mideleg;
  assign T_5868 = pending_interrupts & T_5867;
  assign m_interrupts = T_5866 ? T_5868 : {{63'd0}, 1'h0};
  assign GEN_632 = {{1'd0}, 1'h1};
  assign T_5873 = reg_mstatus_prv < GEN_632;
  assign T_5875 = reg_mstatus_prv == GEN_632;
  assign T_5876 = T_5875 & reg_mstatus_sie;
  assign T_5877 = T_5873 | T_5876;
  assign T_5878 = T_5859 & T_5877;
  assign T_5879 = pending_interrupts & reg_mideleg;
  assign s_interrupts = T_5878 ? T_5879 : {{63'd0}, 1'h0};
  assign all_interrupts = m_interrupts | s_interrupts;
  assign T_5882 = all_interrupts[0];
  assign T_5883 = all_interrupts[1];
  assign T_5884 = all_interrupts[2];
  assign T_5885 = all_interrupts[3];
  assign T_5886 = all_interrupts[4];
  assign T_5887 = all_interrupts[5];
  assign T_5888 = all_interrupts[6];
  assign T_5889 = all_interrupts[7];
  assign T_5890 = all_interrupts[8];
  assign T_5891 = all_interrupts[9];
  assign T_5892 = all_interrupts[10];
  assign T_5893 = all_interrupts[11];
  assign T_5894 = all_interrupts[12];
  assign T_5895 = all_interrupts[13];
  assign T_5896 = all_interrupts[14];
  assign T_5897 = all_interrupts[15];
  assign T_5898 = all_interrupts[16];
  assign T_5899 = all_interrupts[17];
  assign T_5900 = all_interrupts[18];
  assign T_5901 = all_interrupts[19];
  assign T_5902 = all_interrupts[20];
  assign T_5903 = all_interrupts[21];
  assign T_5904 = all_interrupts[22];
  assign T_5905 = all_interrupts[23];
  assign T_5906 = all_interrupts[24];
  assign T_5907 = all_interrupts[25];
  assign T_5908 = all_interrupts[26];
  assign T_5909 = all_interrupts[27];
  assign T_5910 = all_interrupts[28];
  assign T_5911 = all_interrupts[29];
  assign T_5912 = all_interrupts[30];
  assign T_5913 = all_interrupts[31];
  assign T_5914 = all_interrupts[32];
  assign T_5915 = all_interrupts[33];
  assign T_5916 = all_interrupts[34];
  assign T_5917 = all_interrupts[35];
  assign T_5918 = all_interrupts[36];
  assign T_5919 = all_interrupts[37];
  assign T_5920 = all_interrupts[38];
  assign T_5921 = all_interrupts[39];
  assign T_5922 = all_interrupts[40];
  assign T_5923 = all_interrupts[41];
  assign T_5924 = all_interrupts[42];
  assign T_5925 = all_interrupts[43];
  assign T_5926 = all_interrupts[44];
  assign T_5927 = all_interrupts[45];
  assign T_5928 = all_interrupts[46];
  assign T_5929 = all_interrupts[47];
  assign T_5930 = all_interrupts[48];
  assign T_5931 = all_interrupts[49];
  assign T_5932 = all_interrupts[50];
  assign T_5933 = all_interrupts[51];
  assign T_5934 = all_interrupts[52];
  assign T_5935 = all_interrupts[53];
  assign T_5936 = all_interrupts[54];
  assign T_5937 = all_interrupts[55];
  assign T_5938 = all_interrupts[56];
  assign T_5939 = all_interrupts[57];
  assign T_5940 = all_interrupts[58];
  assign T_5941 = all_interrupts[59];
  assign T_5942 = all_interrupts[60];
  assign T_5943 = all_interrupts[61];
  assign T_5944 = all_interrupts[62];
  assign T_6010 = T_5944 ? 6'h3e : 6'h3f;
  assign T_6011 = T_5943 ? 6'h3d : T_6010;
  assign T_6012 = T_5942 ? 6'h3c : T_6011;
  assign T_6013 = T_5941 ? 6'h3b : T_6012;
  assign T_6014 = T_5940 ? 6'h3a : T_6013;
  assign T_6015 = T_5939 ? 6'h39 : T_6014;
  assign T_6016 = T_5938 ? 6'h38 : T_6015;
  assign T_6017 = T_5937 ? 6'h37 : T_6016;
  assign T_6018 = T_5936 ? 6'h36 : T_6017;
  assign T_6019 = T_5935 ? 6'h35 : T_6018;
  assign T_6020 = T_5934 ? 6'h34 : T_6019;
  assign T_6021 = T_5933 ? 6'h33 : T_6020;
  assign T_6022 = T_5932 ? 6'h32 : T_6021;
  assign T_6023 = T_5931 ? 6'h31 : T_6022;
  assign T_6024 = T_5930 ? 6'h30 : T_6023;
  assign T_6025 = T_5929 ? 6'h2f : T_6024;
  assign T_6026 = T_5928 ? 6'h2e : T_6025;
  assign T_6027 = T_5927 ? 6'h2d : T_6026;
  assign T_6028 = T_5926 ? 6'h2c : T_6027;
  assign T_6029 = T_5925 ? 6'h2b : T_6028;
  assign T_6030 = T_5924 ? 6'h2a : T_6029;
  assign T_6031 = T_5923 ? 6'h29 : T_6030;
  assign T_6032 = T_5922 ? 6'h28 : T_6031;
  assign T_6033 = T_5921 ? 6'h27 : T_6032;
  assign T_6034 = T_5920 ? 6'h26 : T_6033;
  assign T_6035 = T_5919 ? 6'h25 : T_6034;
  assign T_6036 = T_5918 ? 6'h24 : T_6035;
  assign T_6037 = T_5917 ? 6'h23 : T_6036;
  assign T_6038 = T_5916 ? 6'h22 : T_6037;
  assign T_6039 = T_5915 ? 6'h21 : T_6038;
  assign T_6040 = T_5914 ? 6'h20 : T_6039;
  assign T_6041 = T_5913 ? {{1'd0}, 5'h1f} : T_6040;
  assign T_6042 = T_5912 ? {{1'd0}, 5'h1e} : T_6041;
  assign T_6043 = T_5911 ? {{1'd0}, 5'h1d} : T_6042;
  assign T_6044 = T_5910 ? {{1'd0}, 5'h1c} : T_6043;
  assign T_6045 = T_5909 ? {{1'd0}, 5'h1b} : T_6044;
  assign T_6046 = T_5908 ? {{1'd0}, 5'h1a} : T_6045;
  assign T_6047 = T_5907 ? {{1'd0}, 5'h19} : T_6046;
  assign T_6048 = T_5906 ? {{1'd0}, 5'h18} : T_6047;
  assign T_6049 = T_5905 ? {{1'd0}, 5'h17} : T_6048;
  assign T_6050 = T_5904 ? {{1'd0}, 5'h16} : T_6049;
  assign T_6051 = T_5903 ? {{1'd0}, 5'h15} : T_6050;
  assign T_6052 = T_5902 ? {{1'd0}, 5'h14} : T_6051;
  assign T_6053 = T_5901 ? {{1'd0}, 5'h13} : T_6052;
  assign T_6054 = T_5900 ? {{1'd0}, 5'h12} : T_6053;
  assign T_6055 = T_5899 ? {{1'd0}, 5'h11} : T_6054;
  assign T_6056 = T_5898 ? {{1'd0}, 5'h10} : T_6055;
  assign T_6057 = T_5897 ? {{2'd0}, 4'hf} : T_6056;
  assign T_6058 = T_5896 ? {{2'd0}, 4'he} : T_6057;
  assign T_6059 = T_5895 ? {{2'd0}, 4'hd} : T_6058;
  assign T_6060 = T_5894 ? {{2'd0}, 4'hc} : T_6059;
  assign T_6061 = T_5893 ? {{2'd0}, 4'hb} : T_6060;
  assign T_6062 = T_5892 ? {{2'd0}, 4'ha} : T_6061;
  assign T_6063 = T_5891 ? {{2'd0}, 4'h9} : T_6062;
  assign T_6064 = T_5890 ? {{2'd0}, 4'h8} : T_6063;
  assign T_6065 = T_5889 ? {{3'd0}, 3'h7} : T_6064;
  assign T_6066 = T_5888 ? {{3'd0}, 3'h6} : T_6065;
  assign T_6067 = T_5887 ? {{3'd0}, 3'h5} : T_6066;
  assign T_6068 = T_5886 ? {{3'd0}, 3'h4} : T_6067;
  assign T_6069 = T_5885 ? {{4'd0}, 2'h3} : T_6068;
  assign T_6070 = T_5884 ? {{4'd0}, 2'h2} : T_6069;
  assign T_6071 = T_5883 ? {{5'd0}, 1'h1} : T_6070;
  assign T_6072 = T_5882 ? {{5'd0}, 1'h0} : T_6071;
  assign GEN_634 = {{58'd0}, T_6072};
  assign T_6073 = 64'h8000000000000000 + GEN_634;
  assign interruptCause = T_6073[63:0];
  assign GEN_635 = {{63'd0}, 1'h0};
  assign T_6075 = all_interrupts != GEN_635;
  assign T_6078 = T_6075 & T_5325;
  assign T_6079 = T_6078 | reg_singleStepped;
  assign T_6084 = reg_dcsr_debugint & T_5859;
  assign GEN_65 = T_6084 ? 1'h1 : T_6079;
  assign GEN_66 = T_6084 ? 64'h800000000000000d : interruptCause;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T_6087 = io_rw_cmd != 3'h0;
  assign T_6089 = system_insn == 1'h0;
  assign cpu_ren = T_6087 & T_6089;
  assign T_6090 = {io_status_sie,io_status_uie};
  assign T_6091 = {io_status_upie,io_status_mie};
  assign T_6092 = {T_6091,io_status_hie};
  assign T_6093 = {T_6092,T_6090};
  assign T_6094 = {io_status_mpie,io_status_hpie};
  assign T_6095 = {T_6094,io_status_spie};
  assign T_6096 = {io_status_mpp,io_status_hpp};
  assign T_6097 = {T_6096,io_status_spp};
  assign T_6098 = {T_6097,T_6095};
  assign T_6099 = {T_6098,T_6093};
  assign T_6100 = {io_status_mprv,io_status_xs};
  assign T_6101 = {T_6100,io_status_fs};
  assign T_6102 = {io_status_vm,io_status_zero1};
  assign T_6103 = {T_6102,io_status_pum};
  assign T_6104 = {T_6103,T_6101};
  assign T_6105 = {io_status_zero3,io_status_sd_rv32};
  assign T_6106 = {T_6105,io_status_zero2};
  assign T_6107 = {io_status_debug,io_status_prv};
  assign T_6108 = {T_6107,io_status_sd};
  assign T_6109 = {T_6108,T_6106};
  assign T_6110 = {T_6109,T_6104};
  assign T_6111 = {T_6110,T_6099};
  assign read_mstatus = T_6111[63:0];
  assign T_6112 = {reg_tdrselect_tdrmode,reg_tdrselect_reserved};
  assign T_6113 = {T_6112,reg_tdrselect_tdrindex};
  assign GEN_0 = GEN_67;
  assign GEN_67 = reg_tdrselect_tdrindex ? reg_bp_1_control_r : reg_bp_0_control_r;
  assign GEN_1 = GEN_68;
  assign GEN_68 = reg_tdrselect_tdrindex ? reg_bp_1_control_w : reg_bp_0_control_w;
  assign T_6128 = {GEN_0,GEN_1};
  assign GEN_2 = GEN_69;
  assign GEN_69 = reg_tdrselect_tdrindex ? reg_bp_1_control_x : reg_bp_0_control_x;
  assign T_6129 = {T_6128,GEN_2};
  assign GEN_3 = GEN_70;
  assign GEN_70 = reg_tdrselect_tdrindex ? reg_bp_1_control_h : reg_bp_0_control_h;
  assign GEN_4 = GEN_71;
  assign GEN_71 = reg_tdrselect_tdrindex ? reg_bp_1_control_s : reg_bp_0_control_s;
  assign T_6130 = {GEN_3,GEN_4};
  assign GEN_5 = GEN_72;
  assign GEN_72 = reg_tdrselect_tdrindex ? reg_bp_1_control_u : reg_bp_0_control_u;
  assign T_6131 = {T_6130,GEN_5};
  assign T_6132 = {T_6131,T_6129};
  assign GEN_6 = GEN_73;
  assign GEN_73 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpaction : reg_bp_0_control_bpaction;
  assign GEN_7 = GEN_74;
  assign GEN_74 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpmatch : reg_bp_0_control_bpmatch;
  assign T_6133 = {GEN_6,GEN_7};
  assign GEN_8 = GEN_75;
  assign GEN_75 = reg_tdrselect_tdrindex ? reg_bp_1_control_m : reg_bp_0_control_m;
  assign T_6134 = {T_6133,GEN_8};
  assign GEN_9 = GEN_76;
  assign GEN_76 = reg_tdrselect_tdrindex ? reg_bp_1_control_tdrtype : reg_bp_0_control_tdrtype;
  assign GEN_10 = GEN_77;
  assign GEN_77 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpamaskmax : reg_bp_0_control_bpamaskmax;
  assign T_6135 = {GEN_9,GEN_10};
  assign GEN_11 = GEN_78;
  assign GEN_78 = reg_tdrselect_tdrindex ? reg_bp_1_control_reserved : reg_bp_0_control_reserved;
  assign T_6136 = {T_6135,GEN_11};
  assign T_6137 = {T_6136,T_6134};
  assign T_6138 = {T_6137,T_6132};
  assign T_6161 = reg_mepc[39];
  assign GEN_636 = {{23'd0}, T_6161};
  assign T_6163 = 24'h0 - GEN_636;
  assign T_6164 = T_6163[23:0];
  assign T_6165 = {T_6164,reg_mepc};
  assign T_6166 = reg_mbadaddr[39];
  assign GEN_637 = {{23'd0}, T_6166};
  assign T_6168 = 24'h0 - GEN_637;
  assign T_6169 = T_6168[23:0];
  assign T_6170 = {T_6169,reg_mbadaddr};
  assign T_6171 = {reg_dcsr_step,reg_dcsr_prv};
  assign T_6172 = {reg_dcsr_zero1,reg_dcsr_halt};
  assign T_6173 = {T_6172,T_6171};
  assign T_6174 = {reg_dcsr_cause,reg_dcsr_debugint};
  assign T_6175 = {reg_dcsr_stopcycle,reg_dcsr_stoptime};
  assign T_6176 = {T_6175,T_6174};
  assign T_6177 = {T_6176,T_6173};
  assign T_6178 = {reg_dcsr_ebreaku,reg_dcsr_zero2};
  assign T_6179 = {reg_dcsr_ebreakh,reg_dcsr_ebreaks};
  assign T_6180 = {T_6179,T_6178};
  assign T_6181 = {reg_dcsr_hwbpcount,reg_dcsr_ebreakm};
  assign T_6182 = {reg_dcsr_xdebugver,reg_dcsr_ndreset};
  assign T_6183 = {T_6182,reg_dcsr_fullreset};
  assign T_6184 = {T_6183,T_6181};
  assign T_6185 = {T_6184,T_6180};
  assign T_6186 = {T_6185,T_6177};
  assign T_6187 = reg_mie & reg_mideleg;
  assign T_6188 = GEN_631 & reg_mideleg;
  assign T_6189_debug = io_status_debug;
  assign T_6189_prv = io_status_prv;
  assign T_6189_sd = io_status_sd;
  assign T_6189_zero3 = io_status_zero3;
  assign T_6189_sd_rv32 = io_status_sd_rv32;
  assign T_6189_zero2 = io_status_zero2;
  assign T_6189_vm = {{4'd0}, 1'h0};
  assign T_6189_zero1 = io_status_zero1;
  assign T_6189_pum = io_status_pum;
  assign T_6189_mprv = 1'h0;
  assign T_6189_xs = io_status_xs;
  assign T_6189_fs = io_status_fs;
  assign T_6189_mpp = {{1'd0}, 1'h0};
  assign T_6189_hpp = {{1'd0}, 1'h0};
  assign T_6189_spp = io_status_spp;
  assign T_6189_mpie = 1'h0;
  assign T_6189_hpie = 1'h0;
  assign T_6189_spie = io_status_spie;
  assign T_6189_upie = io_status_upie;
  assign T_6189_mie = 1'h0;
  assign T_6189_hie = 1'h0;
  assign T_6189_sie = io_status_sie;
  assign T_6189_uie = io_status_uie;
  assign T_6221 = {T_6189_sie,T_6189_uie};
  assign T_6222 = {T_6189_upie,T_6189_mie};
  assign T_6223 = {T_6222,T_6189_hie};
  assign T_6224 = {T_6223,T_6221};
  assign T_6225 = {T_6189_mpie,T_6189_hpie};
  assign T_6226 = {T_6225,T_6189_spie};
  assign T_6227 = {T_6189_mpp,T_6189_hpp};
  assign T_6228 = {T_6227,T_6189_spp};
  assign T_6229 = {T_6228,T_6226};
  assign T_6230 = {T_6229,T_6224};
  assign T_6231 = {T_6189_mprv,T_6189_xs};
  assign T_6232 = {T_6231,T_6189_fs};
  assign T_6233 = {T_6189_vm,T_6189_zero1};
  assign T_6234 = {T_6233,T_6189_pum};
  assign T_6235 = {T_6234,T_6232};
  assign T_6236 = {T_6189_zero3,T_6189_sd_rv32};
  assign T_6237 = {T_6236,T_6189_zero2};
  assign T_6238 = {T_6189_debug,T_6189_prv};
  assign T_6239 = {T_6238,T_6189_sd};
  assign T_6240 = {T_6239,T_6237};
  assign T_6241 = {T_6240,T_6235};
  assign T_6242 = {T_6241,T_6230};
  assign T_6243 = T_6242[63:0];
  assign T_6244 = reg_sbadaddr[39];
  assign GEN_639 = {{23'd0}, T_6244};
  assign T_6246 = 24'h0 - GEN_639;
  assign T_6247 = T_6246[23:0];
  assign T_6248 = {T_6247,reg_sbadaddr};
  assign T_6249 = {reg_sptbr_asid,reg_sptbr_ppn};
  assign T_6250 = reg_sepc[39];
  assign GEN_640 = {{23'd0}, T_6250};
  assign T_6252 = 24'h0 - GEN_640;
  assign T_6253 = T_6252[23:0];
  assign T_6254 = {T_6253,reg_sepc};
  assign T_6255 = reg_stvec[38];
  assign GEN_641 = {{24'd0}, T_6255};
  assign T_6257 = 25'h0 - GEN_641;
  assign T_6258 = T_6257[24:0];
  assign T_6259 = {T_6258,reg_stvec};
  assign GEN_642 = {{1'd0}, 11'h7a0};
  assign T_6265 = io_rw_addr == GEN_642;
  assign GEN_643 = {{1'd0}, 11'h7a1};
  assign T_6267 = io_rw_addr == GEN_643;
  assign GEN_644 = {{1'd0}, 11'h7a2};
  assign T_6269 = io_rw_addr == GEN_644;
  assign T_6271 = io_rw_addr == 12'hf13;
  assign T_6273 = io_rw_addr == 12'hf12;
  assign T_6275 = io_rw_addr == 12'hf11;
  assign T_6277 = io_rw_addr == 12'hf00;
  assign T_6279 = io_rw_addr == 12'hf02;
  assign GEN_645 = {{2'd0}, 10'h310};
  assign T_6281 = io_rw_addr == GEN_645;
  assign GEN_646 = {{1'd0}, 11'h701};
  assign T_6283 = io_rw_addr == GEN_646;
  assign GEN_647 = {{1'd0}, 11'h700};
  assign T_6285 = io_rw_addr == GEN_647;
  assign GEN_648 = {{1'd0}, 11'h702};
  assign T_6287 = io_rw_addr == GEN_648;
  assign T_6289 = io_rw_addr == 12'hf10;
  assign GEN_649 = {{2'd0}, 10'h300};
  assign T_6291 = io_rw_addr == GEN_649;
  assign GEN_650 = {{2'd0}, 10'h305};
  assign T_6293 = io_rw_addr == GEN_650;
  assign GEN_651 = {{2'd0}, 10'h344};
  assign T_6295 = io_rw_addr == GEN_651;
  assign GEN_652 = {{2'd0}, 10'h304};
  assign T_6297 = io_rw_addr == GEN_652;
  assign GEN_653 = {{2'd0}, 10'h303};
  assign T_6299 = io_rw_addr == GEN_653;
  assign GEN_654 = {{2'd0}, 10'h302};
  assign T_6301 = io_rw_addr == GEN_654;
  assign GEN_655 = {{2'd0}, 10'h340};
  assign T_6303 = io_rw_addr == GEN_655;
  assign GEN_656 = {{2'd0}, 10'h341};
  assign T_6305 = io_rw_addr == GEN_656;
  assign GEN_657 = {{2'd0}, 10'h343};
  assign T_6307 = io_rw_addr == GEN_657;
  assign GEN_658 = {{2'd0}, 10'h342};
  assign T_6309 = io_rw_addr == GEN_658;
  assign T_6311 = io_rw_addr == 12'hf14;
  assign GEN_659 = {{1'd0}, 11'h7b0};
  assign T_6313 = io_rw_addr == GEN_659;
  assign GEN_660 = {{1'd0}, 11'h7b1};
  assign T_6315 = io_rw_addr == GEN_660;
  assign GEN_661 = {{1'd0}, 11'h7b2};
  assign T_6317 = io_rw_addr == GEN_661;
  assign GEN_662 = {{3'd0}, 9'h100};
  assign T_6319 = io_rw_addr == GEN_662;
  assign GEN_663 = {{3'd0}, 9'h144};
  assign T_6321 = io_rw_addr == GEN_663;
  assign GEN_664 = {{3'd0}, 9'h104};
  assign T_6323 = io_rw_addr == GEN_664;
  assign GEN_665 = {{3'd0}, 9'h140};
  assign T_6325 = io_rw_addr == GEN_665;
  assign GEN_666 = {{3'd0}, 9'h142};
  assign T_6327 = io_rw_addr == GEN_666;
  assign GEN_667 = {{3'd0}, 9'h143};
  assign T_6329 = io_rw_addr == GEN_667;
  assign GEN_668 = {{3'd0}, 9'h180};
  assign T_6331 = io_rw_addr == GEN_668;
  assign GEN_669 = {{3'd0}, 9'h141};
  assign T_6333 = io_rw_addr == GEN_669;
  assign GEN_670 = {{3'd0}, 9'h105};
  assign T_6335 = io_rw_addr == GEN_670;
  assign GEN_671 = {{2'd0}, 10'h311};
  assign T_6337 = io_rw_addr == GEN_671;
  assign GEN_672 = {{1'd0}, 11'h705};
  assign T_6339 = io_rw_addr == GEN_672;
  assign GEN_673 = {{1'd0}, 11'h704};
  assign T_6341 = io_rw_addr == GEN_673;
  assign GEN_674 = {{1'd0}, 11'h706};
  assign T_6343 = io_rw_addr == GEN_674;
  assign T_6344 = T_6265 | T_6267;
  assign T_6345 = T_6344 | T_6269;
  assign T_6346 = T_6345 | T_6271;
  assign T_6347 = T_6346 | T_6273;
  assign T_6348 = T_6347 | T_6275;
  assign T_6349 = T_6348 | T_6277;
  assign T_6350 = T_6349 | T_6279;
  assign T_6351 = T_6350 | T_6281;
  assign T_6352 = T_6351 | T_6283;
  assign T_6353 = T_6352 | T_6285;
  assign T_6354 = T_6353 | T_6287;
  assign T_6355 = T_6354 | T_6289;
  assign T_6356 = T_6355 | T_6291;
  assign T_6357 = T_6356 | T_6293;
  assign T_6358 = T_6357 | T_6295;
  assign T_6359 = T_6358 | T_6297;
  assign T_6360 = T_6359 | T_6299;
  assign T_6361 = T_6360 | T_6301;
  assign T_6362 = T_6361 | T_6303;
  assign T_6363 = T_6362 | T_6305;
  assign T_6364 = T_6363 | T_6307;
  assign T_6365 = T_6364 | T_6309;
  assign T_6366 = T_6365 | T_6311;
  assign T_6367 = T_6366 | T_6313;
  assign T_6368 = T_6367 | T_6315;
  assign T_6369 = T_6368 | T_6317;
  assign T_6370 = T_6369 | T_6319;
  assign T_6371 = T_6370 | T_6321;
  assign T_6372 = T_6371 | T_6323;
  assign T_6373 = T_6372 | T_6325;
  assign T_6374 = T_6373 | T_6327;
  assign T_6375 = T_6374 | T_6329;
  assign T_6376 = T_6375 | T_6331;
  assign T_6377 = T_6376 | T_6333;
  assign T_6378 = T_6377 | T_6335;
  assign T_6379 = T_6378 | T_6337;
  assign T_6380 = T_6379 | T_6339;
  assign T_6381 = T_6380 | T_6341;
  assign addr_valid = T_6381 | T_6343;
  assign T_6383 = io_rw_addr[5];
  assign T_6384 = io_rw_addr[6:5];
  assign T_6385 = ~ T_6384;
  assign GEN_675 = {{1'd0}, 1'h0};
  assign T_6387 = T_6385 == GEN_675;
  assign T_6388 = io_rw_addr[9:8];
  assign csr_addr_priv = {T_6387,T_6388};
  assign T_6389 = {reg_debug,reg_mstatus_prv};
  assign priv_sufficient = T_6389 >= csr_addr_priv;
  assign T_6390 = io_rw_addr[11:10];
  assign T_6391 = ~ T_6390;
  assign read_only = T_6391 == GEN_675;
  assign T_6393 = io_rw_cmd != 3'h5;
  assign T_6394 = cpu_ren & T_6393;
  assign cpu_wen = T_6394 & priv_sufficient;
  assign T_6396 = read_only == 1'h0;
  assign wen = cpu_wen & T_6396;
  assign T_6397 = io_rw_cmd == 3'h2;
  assign T_6398 = io_rw_cmd == 3'h3;
  assign T_6399 = T_6397 | T_6398;
  assign T_6401 = T_6399 ? io_rw_rdata : {{63'd0}, 1'h0};
  assign T_6402 = io_rw_cmd != 3'h3;
  assign T_6404 = T_6402 ? io_rw_wdata : {{63'd0}, 1'h0};
  assign T_6405 = T_6401 | T_6404;
  assign T_6408 = T_6398 ? io_rw_wdata : {{63'd0}, 1'h0};
  assign T_6409 = ~ T_6408;
  assign wdata = T_6405 & T_6409;
  assign do_system_insn = priv_sufficient & system_insn;
  assign T_6411 = io_rw_addr[2:0];
  assign GEN_677 = {{7'd0}, 1'h1};
  assign opcode = GEN_677 << T_6411;
  assign T_6412 = opcode[0];
  assign insn_call = do_system_insn & T_6412;
  assign T_6413 = opcode[1];
  assign insn_break = do_system_insn & T_6413;
  assign T_6414 = opcode[2];
  assign insn_ret = do_system_insn & T_6414;
  assign T_6415 = opcode[4];
  assign insn_sfence_vm = do_system_insn & T_6415;
  assign T_6416 = opcode[5];
  assign insn_wfi = do_system_insn & T_6416;
  assign T_6417 = cpu_wen & read_only;
  assign T_6419 = priv_sufficient == 1'h0;
  assign T_6421 = addr_valid == 1'h0;
  assign T_6422 = T_6419 | T_6421;
  assign T_6429 = cpu_ren & T_6422;
  assign T_6430 = T_6417 | T_6429;
  assign T_6433 = system_insn & T_6419;
  assign T_6434 = T_6430 | T_6433;
  assign T_6435 = T_6434 | insn_call;
  assign T_6436 = T_6435 | insn_break;
  assign GEN_79 = insn_wfi ? 1'h1 : reg_wfi;
  assign GEN_679 = {{12'd0}, 1'h0};
  assign T_6439 = read_mip != GEN_679;
  assign GEN_80 = T_6439 ? 1'h0 : GEN_79;
  assign T_6442 = io_csr_xcpt == 1'h0;
  assign GEN_680 = {{2'd0}, reg_mstatus_prv};
  assign T_6444 = GEN_680 + 4'h8;
  assign T_6445 = T_6444[3:0];
  assign T_6448 = insn_break ? 2'h3 : 2'h2;
  assign T_6449 = insn_call ? T_6445 : {{2'd0}, T_6448};
  assign cause = T_6442 ? io_cause : {{60'd0}, T_6449};
  assign cause_lsbs = cause[5:0];
  assign T_6450 = cause[63];
  assign GEN_681 = {{2'd0}, 4'hd};
  assign T_6452 = cause_lsbs == GEN_681;
  assign causeIsDebugInt = T_6450 & T_6452;
  assign GEN_682 = {{62'd0}, 2'h3};
  assign T_6454 = cause == GEN_682;
  assign T_6455 = {reg_dcsr_ebreaks,reg_dcsr_ebreaku};
  assign T_6456 = {reg_dcsr_ebreakm,reg_dcsr_ebreakh};
  assign T_6457 = {T_6456,T_6455};
  assign T_6458 = T_6457 >> reg_mstatus_prv;
  assign T_6459 = T_6458[0];
  assign causeIsDebugBreak = T_6454 & T_6459;
  assign T_6461 = reg_singleStepped | causeIsDebugInt;
  assign T_6462 = T_6461 | causeIsDebugBreak;
  assign T_6463 = T_6462 | reg_debug;
  assign T_6469 = reg_mideleg >> cause_lsbs;
  assign T_6470 = T_6469[0];
  assign T_6471 = reg_medeleg >> cause_lsbs;
  assign T_6472 = T_6471[0];
  assign T_6473 = T_6450 ? T_6470 : T_6472;
  assign delegate = T_5861 & T_6473;
  assign debugTVec = reg_debug ? 12'h808 : 12'h800;
  assign T_6477 = {T_6255,reg_stvec};
  assign T_6478 = delegate ? T_6477 : {{8'd0}, reg_mtvec};
  assign tvec = T_6463 ? {{28'd0}, debugTVec} : T_6478;
  assign T_6480 = csr_addr_priv[1];
  assign T_6482 = T_6480 == 1'h0;
  assign T_6484 = T_6482 ? reg_sepc : reg_mepc;
  assign epc = T_6383 ? reg_dpc : T_6484;
  assign T_6485 = exception ? tvec : epc;
  assign T_6488 = reg_dcsr_step & T_5859;
  assign T_6489 = ~ io_status_fs;
  assign T_6491 = T_6489 == GEN_675;
  assign T_6492 = ~ io_status_xs;
  assign T_6494 = T_6492 == GEN_675;
  assign T_6495 = T_6491 | T_6494;
  assign T_6496 = ~ io_pc;
  assign GEN_685 = {{38'd0}, 2'h3};
  assign T_6498 = T_6496 | GEN_685;
  assign T_6499 = ~ T_6498;
  assign T_6500 = read_mstatus >> reg_mstatus_prv;
  assign T_6501 = T_6500[0];
  assign T_6506 = causeIsDebugInt ? 2'h3 : {{1'd0}, 1'h1};
  assign T_6507 = reg_singleStepped ? 3'h4 : {{1'd0}, T_6506};
  assign GEN_81 = T_6463 ? 1'h1 : reg_debug;
  assign GEN_82 = T_6463 ? T_6499 : reg_dpc;
  assign GEN_83 = T_6463 ? T_6507 : reg_dcsr_cause;
  assign GEN_84 = T_6463 ? reg_mstatus_prv : reg_dcsr_prv;
  assign T_6509 = T_6463 == 1'h0;
  assign T_6510 = T_6509 & delegate;
  assign GEN_85 = T_6510 ? T_6499 : reg_sepc;
  assign GEN_86 = T_6510 ? cause : reg_scause;
  assign GEN_87 = T_6510 ? io_badaddr : reg_sbadaddr;
  assign GEN_88 = T_6510 ? T_6501 : reg_mstatus_spie;
  assign GEN_89 = T_6510 ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp};
  assign GEN_90 = T_6510 ? 1'h0 : reg_mstatus_sie;
  assign GEN_91 = T_6510 ? {{1'd0}, 1'h1} : reg_mstatus_prv;
  assign T_6516 = delegate == 1'h0;
  assign T_6517 = T_6509 & T_6516;
  assign GEN_92 = T_6517 ? T_6499 : reg_mepc;
  assign GEN_93 = T_6517 ? cause : reg_mcause;
  assign GEN_94 = T_6517 ? io_badaddr : reg_mbadaddr;
  assign GEN_95 = T_6517 ? T_6501 : reg_mstatus_mpie;
  assign GEN_96 = T_6517 ? reg_mstatus_prv : reg_mstatus_mpp;
  assign GEN_97 = T_6517 ? 1'h0 : reg_mstatus_mie;
  assign GEN_98 = T_6517 ? 2'h3 : GEN_91;
  assign GEN_99 = exception ? GEN_81 : reg_debug;
  assign GEN_100 = exception ? GEN_82 : reg_dpc;
  assign GEN_101 = exception ? GEN_83 : reg_dcsr_cause;
  assign GEN_102 = exception ? GEN_84 : reg_dcsr_prv;
  assign GEN_103 = exception ? GEN_85 : reg_sepc;
  assign GEN_104 = exception ? GEN_86 : reg_scause;
  assign GEN_105 = exception ? GEN_87 : reg_sbadaddr;
  assign GEN_106 = exception ? GEN_88 : reg_mstatus_spie;
  assign GEN_107 = exception ? GEN_89 : {{1'd0}, reg_mstatus_spp};
  assign GEN_108 = exception ? GEN_90 : reg_mstatus_sie;
  assign GEN_109 = exception ? GEN_98 : reg_mstatus_prv;
  assign GEN_110 = exception ? GEN_92 : reg_mepc;
  assign GEN_111 = exception ? GEN_93 : reg_mcause;
  assign GEN_112 = exception ? GEN_94 : reg_mbadaddr;
  assign GEN_113 = exception ? GEN_95 : reg_mstatus_mpie;
  assign GEN_114 = exception ? GEN_96 : reg_mstatus_mpp;
  assign GEN_115 = exception ? GEN_97 : reg_mstatus_mie;
  assign GEN_116 = reg_mstatus_spp ? reg_mstatus_spie : GEN_108;
  assign GEN_117 = T_6482 ? GEN_116 : GEN_108;
  assign GEN_118 = T_6482 ? 1'h0 : GEN_106;
  assign GEN_119 = T_6482 ? {{1'd0}, 1'h0} : GEN_107;
  assign GEN_120 = T_6482 ? {{1'd0}, reg_mstatus_spp} : GEN_109;
  assign T_6529 = T_6482 == 1'h0;
  assign T_6530 = T_6529 & T_6383;
  assign GEN_121 = T_6530 ? reg_dcsr_prv : GEN_120;
  assign GEN_122 = T_6530 ? 1'h0 : GEN_99;
  assign T_6535 = T_6383 == 1'h0;
  assign T_6536 = T_6529 & T_6535;
  assign T_6537 = reg_mstatus_mpp[1];
  assign GEN_123 = T_6537 ? reg_mstatus_mpie : GEN_115;
  assign T_6539 = reg_mstatus_mpp[0];
  assign T_6542 = T_6537 == 1'h0;
  assign T_6543 = T_6542 & T_6539;
  assign GEN_124 = T_6543 ? reg_mstatus_mpie : GEN_117;
  assign GEN_125 = T_6536 ? GEN_123 : GEN_115;
  assign GEN_126 = T_6536 ? GEN_124 : GEN_117;
  assign GEN_127 = T_6536 ? 1'h0 : GEN_113;
  assign GEN_128 = T_6536 ? {{1'd0}, 1'h0} : GEN_114;
  assign GEN_129 = T_6536 ? reg_mstatus_mpp : GEN_121;
  assign GEN_130 = insn_ret ? GEN_126 : GEN_108;
  assign GEN_131 = insn_ret ? GEN_118 : GEN_106;
  assign GEN_132 = insn_ret ? GEN_119 : GEN_107;
  assign GEN_133 = insn_ret ? GEN_129 : GEN_109;
  assign GEN_134 = insn_ret ? GEN_122 : GEN_99;
  assign GEN_135 = insn_ret ? GEN_125 : GEN_115;
  assign GEN_136 = insn_ret ? GEN_127 : GEN_113;
  assign GEN_137 = insn_ret ? GEN_128 : GEN_114;
  assign T_6548 = {1'h0,io_csr_xcpt};
  assign GEN_686 = {{1'd0}, io_exception};
  assign T_6549 = GEN_686 + T_6548;
  assign T_6550 = T_6549[1:0];
  assign T_6551 = {1'h0,T_6550};
  assign GEN_687 = {{2'd0}, insn_ret};
  assign T_6552 = GEN_687 + T_6551;
  assign T_6553 = T_6552[2:0];
  assign GEN_688 = {{2'd0}, 1'h1};
  assign T_6555 = T_6553 <= GEN_688;
  assign T_6556 = T_6555 | reset;
  assign T_6558 = T_6556 == 1'h0;
  assign T_6560 = T_6265 ? T_6113 : {{63'd0}, 1'h0};
  assign T_6562 = T_6267 ? T_6138 : {{63'd0}, 1'h0};
  assign GEN_12 = GEN_138;
  assign GEN_138 = reg_tdrselect_tdrindex ? reg_bp_1_address : reg_bp_0_address;
  assign T_6564 = T_6269 ? GEN_12 : {{38'd0}, 1'h0};
  assign T_6572 = T_6277 ? reg_cycle : {{63'd0}, 1'h0};
  assign T_6574 = T_6279 ? T_5816 : {{63'd0}, 1'h0};
  assign T_6584 = T_6289 ? 64'h8000000000041101 : {{63'd0}, 1'h0};
  assign T_6586 = T_6291 ? read_mstatus : {{63'd0}, 1'h0};
  assign T_6588 = T_6293 ? reg_mtvec : {{31'd0}, 1'h0};
  assign T_6590 = T_6295 ? read_mip : {{12'd0}, 1'h0};
  assign T_6592 = T_6297 ? reg_mie : {{63'd0}, 1'h0};
  assign T_6594 = T_6299 ? reg_mideleg : {{63'd0}, 1'h0};
  assign T_6596 = T_6301 ? reg_medeleg : {{63'd0}, 1'h0};
  assign T_6598 = T_6303 ? reg_mscratch : {{63'd0}, 1'h0};
  assign T_6600 = T_6305 ? T_6165 : {{63'd0}, 1'h0};
  assign T_6602 = T_6307 ? T_6170 : {{63'd0}, 1'h0};
  assign T_6604 = T_6309 ? reg_mcause : {{63'd0}, 1'h0};
  assign T_6606 = T_6311 ? io_prci_id : 1'h0;
  assign T_6608 = T_6313 ? T_6186 : {{31'd0}, 1'h0};
  assign T_6610 = T_6315 ? reg_dpc : {{39'd0}, 1'h0};
  assign T_6612 = T_6317 ? reg_dscratch : {{63'd0}, 1'h0};
  assign T_6614 = T_6319 ? T_6243 : {{63'd0}, 1'h0};
  assign T_6616 = T_6321 ? T_6188 : {{63'd0}, 1'h0};
  assign T_6618 = T_6323 ? T_6187 : {{63'd0}, 1'h0};
  assign T_6620 = T_6325 ? reg_sscratch : {{63'd0}, 1'h0};
  assign T_6622 = T_6327 ? reg_scause : {{63'd0}, 1'h0};
  assign T_6624 = T_6329 ? T_6248 : {{63'd0}, 1'h0};
  assign T_6626 = T_6331 ? T_6249 : {{44'd0}, 1'h0};
  assign T_6628 = T_6333 ? T_6254 : {{63'd0}, 1'h0};
  assign T_6630 = T_6335 ? T_6259 : {{63'd0}, 1'h0};
  assign T_6640 = T_6560 | T_6562;
  assign GEN_689 = {{25'd0}, T_6564};
  assign T_6641 = T_6640 | GEN_689;
  assign T_6642 = T_6641 | GEN_635;
  assign T_6643 = T_6642 | GEN_635;
  assign T_6644 = T_6643 | GEN_635;
  assign T_6645 = T_6644 | T_6572;
  assign T_6646 = T_6645 | T_6574;
  assign T_6647 = T_6646 | GEN_635;
  assign T_6648 = T_6647 | GEN_635;
  assign T_6649 = T_6648 | GEN_635;
  assign T_6650 = T_6649 | GEN_635;
  assign T_6651 = T_6650 | T_6584;
  assign T_6652 = T_6651 | T_6586;
  assign GEN_697 = {{32'd0}, T_6588};
  assign T_6653 = T_6652 | GEN_697;
  assign GEN_698 = {{51'd0}, T_6590};
  assign T_6654 = T_6653 | GEN_698;
  assign T_6655 = T_6654 | T_6592;
  assign T_6656 = T_6655 | T_6594;
  assign T_6657 = T_6656 | T_6596;
  assign T_6658 = T_6657 | T_6598;
  assign T_6659 = T_6658 | T_6600;
  assign T_6660 = T_6659 | T_6602;
  assign T_6661 = T_6660 | T_6604;
  assign GEN_699 = {{63'd0}, T_6606};
  assign T_6662 = T_6661 | GEN_699;
  assign GEN_700 = {{32'd0}, T_6608};
  assign T_6663 = T_6662 | GEN_700;
  assign GEN_701 = {{24'd0}, T_6610};
  assign T_6664 = T_6663 | GEN_701;
  assign T_6665 = T_6664 | T_6612;
  assign T_6666 = T_6665 | T_6614;
  assign T_6667 = T_6666 | T_6616;
  assign T_6668 = T_6667 | T_6618;
  assign T_6669 = T_6668 | T_6620;
  assign T_6670 = T_6669 | T_6622;
  assign T_6671 = T_6670 | T_6624;
  assign GEN_702 = {{19'd0}, T_6626};
  assign T_6672 = T_6671 | GEN_702;
  assign T_6673 = T_6672 | T_6628;
  assign T_6674 = T_6673 | T_6630;
  assign T_6675 = T_6674 | GEN_635;
  assign T_6676 = T_6675 | GEN_635;
  assign T_6677 = T_6676 | GEN_635;
  assign T_6678 = T_6677 | GEN_635;
  assign T_6679 = T_6678;
  assign T_6680 = reg_fflags | io_fcsr_flags_bits;
  assign GEN_139 = io_fcsr_flags_valid ? T_6680 : reg_fflags;
  assign supportedModes_0 = 2'h3;
  assign supportedModes_1 = {{1'd0}, 1'h0};
  assign supportedModes_2 = {{1'd0}, 1'h1};
  assign T_6738_debug = T_6786;
  assign T_6738_prv = T_6785;
  assign T_6738_sd = T_6784;
  assign T_6738_zero3 = T_6783;
  assign T_6738_sd_rv32 = T_6782;
  assign T_6738_zero2 = T_6781;
  assign T_6738_vm = T_6780;
  assign T_6738_zero1 = T_6779;
  assign T_6738_pum = T_6778;
  assign T_6738_mprv = T_6777;
  assign T_6738_xs = T_6776;
  assign T_6738_fs = T_6775;
  assign T_6738_mpp = T_6774;
  assign T_6738_hpp = T_6773;
  assign T_6738_spp = T_6772;
  assign T_6738_mpie = T_6771;
  assign T_6738_hpie = T_6770;
  assign T_6738_spie = T_6769;
  assign T_6738_upie = T_6768;
  assign T_6738_mie = T_6767;
  assign T_6738_hie = T_6766;
  assign T_6738_sie = T_6765;
  assign T_6738_uie = T_6764;
  assign T_6763 = {{3'd0}, wdata};
  assign T_6764 = T_6763[0];
  assign T_6765 = T_6763[1];
  assign T_6766 = T_6763[2];
  assign T_6767 = T_6763[3];
  assign T_6768 = T_6763[4];
  assign T_6769 = T_6763[5];
  assign T_6770 = T_6763[6];
  assign T_6771 = T_6763[7];
  assign T_6772 = T_6763[8];
  assign T_6773 = T_6763[10:9];
  assign T_6774 = T_6763[12:11];
  assign T_6775 = T_6763[14:13];
  assign T_6776 = T_6763[16:15];
  assign T_6777 = T_6763[17];
  assign T_6778 = T_6763[18];
  assign T_6779 = T_6763[23:19];
  assign T_6780 = T_6763[28:24];
  assign T_6781 = T_6763[30:29];
  assign T_6782 = T_6763[31];
  assign T_6783 = T_6763[62:32];
  assign T_6784 = T_6763[63];
  assign T_6785 = T_6763[65:64];
  assign T_6786 = T_6763[66];
  assign T_6787 = supportedModes_0 == T_6738_mpp;
  assign T_6788 = supportedModes_1 == T_6738_mpp;
  assign T_6789 = supportedModes_2 == T_6738_mpp;
  assign T_6792 = T_6787 | T_6788;
  assign T_6793 = T_6792 | T_6789;
  assign GEN_140 = T_6793 ? T_6738_mpp : GEN_137;
  assign GEN_707 = {{4'd0}, 1'h0};
  assign T_6795 = T_6738_vm == GEN_707;
  assign GEN_141 = T_6795 ? {{4'd0}, 1'h0} : reg_mstatus_vm;
  assign GEN_708 = {{1'd0}, 4'h9};
  assign T_6798 = T_6738_vm == GEN_708;
  assign GEN_142 = T_6798 ? {{1'd0}, 4'h9} : GEN_141;
  assign T_6801 = T_6738_fs != GEN_675;
  assign GEN_710 = {{1'd0}, T_6801};
  assign T_6803 = 2'h0 - GEN_710;
  assign T_6804 = T_6803[1:0];
  assign GEN_167 = T_6291 ? T_6738_mie : GEN_135;
  assign GEN_168 = T_6291 ? T_6738_mpie : GEN_136;
  assign GEN_169 = T_6291 ? T_6738_mprv : reg_mstatus_mprv;
  assign GEN_170 = T_6291 ? GEN_140 : GEN_137;
  assign GEN_171 = T_6291 ? T_6738_pum : reg_mstatus_pum;
  assign GEN_172 = T_6291 ? {{1'd0}, T_6738_spp} : GEN_132;
  assign GEN_173 = T_6291 ? T_6738_spie : GEN_131;
  assign GEN_174 = T_6291 ? T_6738_sie : GEN_130;
  assign GEN_175 = T_6291 ? GEN_142 : reg_mstatus_vm;
  assign GEN_176 = T_6291 ? T_6804 : reg_mstatus_fs;
  assign T_6833_rocc = T_6859;
  assign T_6833_meip = T_6858;
  assign T_6833_heip = T_6857;
  assign T_6833_seip = T_6856;
  assign T_6833_ueip = T_6855;
  assign T_6833_mtip = T_6854;
  assign T_6833_htip = T_6853;
  assign T_6833_stip = T_6852;
  assign T_6833_utip = T_6851;
  assign T_6833_msip = T_6850;
  assign T_6833_hsip = T_6849;
  assign T_6833_ssip = T_6848;
  assign T_6833_usip = T_6847;
  assign T_6847 = wdata[0];
  assign T_6848 = wdata[1];
  assign T_6849 = wdata[2];
  assign T_6850 = wdata[3];
  assign T_6851 = wdata[4];
  assign T_6852 = wdata[5];
  assign T_6853 = wdata[6];
  assign T_6854 = wdata[7];
  assign T_6855 = wdata[8];
  assign T_6856 = wdata[9];
  assign T_6857 = wdata[10];
  assign T_6858 = wdata[11];
  assign T_6859 = wdata[12];
  assign GEN_190 = T_6295 ? T_6833_ssip : reg_mip_ssip;
  assign GEN_191 = T_6295 ? T_6833_stip : reg_mip_stip;
  assign GEN_711 = {{51'd0}, supported_interrupts};
  assign T_6860 = wdata & GEN_711;
  assign GEN_192 = T_6297 ? T_6860 : reg_mie;
  assign T_6861 = ~ wdata;
  assign T_6863 = T_6861 | GEN_682;
  assign T_6864 = ~ T_6863;
  assign GEN_193 = T_6305 ? T_6864 : {{24'd0}, GEN_110};
  assign GEN_194 = T_6303 ? wdata : reg_mscratch;
  assign T_6865 = wdata[63:2];
  assign GEN_713 = {{2'd0}, T_6865};
  assign T_6866 = GEN_713 << 2;
  assign GEN_195 = T_6293 ? T_6866 : {{32'd0}, reg_mtvec};
  assign T_6868 = wdata & 64'h800000000000001f;
  assign GEN_196 = T_6309 ? T_6868 : GEN_111;
  assign T_6869 = wdata[39:0];
  assign GEN_197 = T_6307 ? T_6869 : GEN_112;
  assign T_6906_xdebugver = T_6940;
  assign T_6906_ndreset = T_6939;
  assign T_6906_fullreset = T_6938;
  assign T_6906_hwbpcount = T_6937;
  assign T_6906_ebreakm = T_6936;
  assign T_6906_ebreakh = T_6935;
  assign T_6906_ebreaks = T_6934;
  assign T_6906_ebreaku = T_6859;
  assign T_6906_zero2 = T_6858;
  assign T_6906_stopcycle = T_6857;
  assign T_6906_stoptime = T_6856;
  assign T_6906_cause = T_6929;
  assign T_6906_debugint = T_6852;
  assign T_6906_zero1 = T_6851;
  assign T_6906_halt = T_6850;
  assign T_6906_step = T_6849;
  assign T_6906_prv = T_6924;
  assign T_6924 = wdata[1:0];
  assign T_6929 = wdata[8:6];
  assign T_6934 = wdata[13];
  assign T_6935 = wdata[14];
  assign T_6936 = wdata[15];
  assign T_6937 = wdata[27:16];
  assign T_6938 = wdata[28];
  assign T_6939 = wdata[29];
  assign T_6940 = wdata[31:30];
  assign GEN_215 = T_6313 ? T_6906_halt : reg_dcsr_halt;
  assign GEN_216 = T_6313 ? T_6906_step : reg_dcsr_step;
  assign GEN_217 = T_6313 ? T_6906_ebreakm : reg_dcsr_ebreakm;
  assign GEN_218 = T_6313 ? T_6906_ebreaks : reg_dcsr_ebreaks;
  assign GEN_219 = T_6313 ? T_6906_ebreaku : reg_dcsr_ebreaku;
  assign GEN_220 = T_6313 ? T_6906_prv : GEN_102;
  assign GEN_221 = T_6315 ? T_6864 : {{24'd0}, GEN_100};
  assign GEN_222 = T_6317 ? wdata : reg_dscratch;
  assign T_6993_debug = T_7041;
  assign T_6993_prv = T_7040;
  assign T_6993_sd = T_7039;
  assign T_6993_zero3 = T_7038;
  assign T_6993_sd_rv32 = T_7037;
  assign T_6993_zero2 = T_7036;
  assign T_6993_vm = T_7035;
  assign T_6993_zero1 = T_7034;
  assign T_6993_pum = T_7033;
  assign T_6993_mprv = T_7032;
  assign T_6993_xs = T_7031;
  assign T_6993_fs = T_7030;
  assign T_6993_mpp = T_7029;
  assign T_6993_hpp = T_7028;
  assign T_6993_spp = T_7027;
  assign T_6993_mpie = T_7026;
  assign T_6993_hpie = T_7025;
  assign T_6993_spie = T_7024;
  assign T_6993_upie = T_7023;
  assign T_6993_mie = T_7022;
  assign T_6993_hie = T_7021;
  assign T_6993_sie = T_7020;
  assign T_6993_uie = T_7019;
  assign T_7018 = {{3'd0}, wdata};
  assign T_7019 = T_7018[0];
  assign T_7020 = T_7018[1];
  assign T_7021 = T_7018[2];
  assign T_7022 = T_7018[3];
  assign T_7023 = T_7018[4];
  assign T_7024 = T_7018[5];
  assign T_7025 = T_7018[6];
  assign T_7026 = T_7018[7];
  assign T_7027 = T_7018[8];
  assign T_7028 = T_7018[10:9];
  assign T_7029 = T_7018[12:11];
  assign T_7030 = T_7018[14:13];
  assign T_7031 = T_7018[16:15];
  assign T_7032 = T_7018[17];
  assign T_7033 = T_7018[18];
  assign T_7034 = T_7018[23:19];
  assign T_7035 = T_7018[28:24];
  assign T_7036 = T_7018[30:29];
  assign T_7037 = T_7018[31];
  assign T_7038 = T_7018[62:32];
  assign T_7039 = T_7018[63];
  assign T_7040 = T_7018[65:64];
  assign T_7041 = T_7018[66];
  assign T_7043 = T_6993_fs != GEN_675;
  assign GEN_716 = {{1'd0}, T_7043};
  assign T_7045 = 2'h0 - GEN_716;
  assign T_7046 = T_7045[1:0];
  assign GEN_247 = T_6319 ? T_6993_sie : GEN_174;
  assign GEN_248 = T_6319 ? T_6993_spie : GEN_173;
  assign GEN_249 = T_6319 ? {{1'd0}, T_6993_spp} : GEN_172;
  assign GEN_250 = T_6319 ? T_6993_pum : GEN_171;
  assign GEN_251 = T_6319 ? T_7046 : GEN_176;
  assign T_7075_rocc = T_6859;
  assign T_7075_meip = T_6858;
  assign T_7075_heip = T_6857;
  assign T_7075_seip = T_6856;
  assign T_7075_ueip = T_6855;
  assign T_7075_mtip = T_6854;
  assign T_7075_htip = T_6853;
  assign T_7075_stip = T_6852;
  assign T_7075_utip = T_6851;
  assign T_7075_msip = T_6850;
  assign T_7075_hsip = T_6849;
  assign T_7075_ssip = T_6848;
  assign T_7075_usip = T_6847;
  assign GEN_265 = T_6321 ? T_7075_ssip : GEN_190;
  assign T_7103 = reg_mie & T_5867;
  assign T_7104 = wdata & reg_mideleg;
  assign T_7105 = T_7103 | T_7104;
  assign GEN_266 = T_6323 ? T_7105 : GEN_192;
  assign GEN_267 = T_6325 ? wdata : reg_sscratch;
  assign T_7106 = wdata[19:0];
  assign GEN_268 = T_6331 ? {{18'd0}, T_7106} : reg_sptbr_ppn;
  assign GEN_269 = T_6333 ? T_6866 : {{24'd0}, GEN_103};
  assign GEN_270 = T_6335 ? T_6866 : {{25'd0}, reg_stvec};
  assign GEN_271 = T_6327 ? T_6868 : GEN_104;
  assign GEN_272 = T_6329 ? T_6869 : GEN_105;
  assign GEN_719 = {{51'd0}, delegable_interrupts};
  assign T_7114 = wdata & GEN_719;
  assign GEN_273 = T_6299 ? T_7114 : reg_mideleg;
  assign GEN_720 = {{55'd0}, 9'h1ab};
  assign T_7115 = wdata & GEN_720;
  assign GEN_274 = T_6301 ? T_7115 : reg_medeleg;
  assign T_7124_tdrmode = T_7130;
  assign T_7124_reserved = T_7129;
  assign T_7124_tdrindex = T_6847;
  assign T_7129 = wdata[62:1];
  assign T_7130 = wdata[63];
  assign GEN_275 = T_6265 ? T_7124_tdrindex : reg_tdrselect_tdrindex;
  assign T_7131 = reg_tdrselect_tdrmode | reg_debug;
  assign T_7158_tdrtype = T_7182;
  assign T_7158_bpamaskmax = T_7181;
  assign T_7158_reserved = T_7180;
  assign T_7158_bpaction = T_7179;
  assign T_7158_bpmatch = T_7178;
  assign T_7158_m = T_6853;
  assign T_7158_h = T_6852;
  assign T_7158_s = T_6851;
  assign T_7158_u = T_6850;
  assign T_7158_r = T_6849;
  assign T_7158_w = T_6848;
  assign T_7158_x = T_6847;
  assign T_7178 = wdata[10:7];
  assign T_7179 = wdata[18:11];
  assign T_7180 = wdata[54:19];
  assign T_7181 = wdata[59:55];
  assign T_7182 = wdata[63:60];
  assign GEN_13 = T_7158_tdrtype;
  assign GEN_14 = T_7158_bpamaskmax;
  assign GEN_15 = T_7158_reserved;
  assign GEN_16 = T_7158_bpaction;
  assign GEN_17 = T_7158_bpmatch;
  assign GEN_284 = 1'h0 == reg_tdrselect_tdrindex ? GEN_17 : reg_bp_0_control_bpmatch;
  assign GEN_18 = T_7158_m;
  assign GEN_286 = 1'h0 == reg_tdrselect_tdrindex ? GEN_18 : reg_bp_0_control_m;
  assign GEN_19 = T_7158_h;
  assign GEN_20 = T_7158_s;
  assign GEN_290 = 1'h0 == reg_tdrselect_tdrindex ? GEN_20 : reg_bp_0_control_s;
  assign GEN_21 = T_7158_u;
  assign GEN_292 = 1'h0 == reg_tdrselect_tdrindex ? GEN_21 : reg_bp_0_control_u;
  assign GEN_22 = T_7158_r;
  assign GEN_294 = 1'h0 == reg_tdrselect_tdrindex ? GEN_22 : reg_bp_0_control_r;
  assign GEN_23 = T_7158_w;
  assign GEN_296 = 1'h0 == reg_tdrselect_tdrindex ? GEN_23 : reg_bp_0_control_w;
  assign GEN_24 = T_7158_x;
  assign GEN_298 = 1'h0 == reg_tdrselect_tdrindex ? GEN_24 : reg_bp_0_control_x;
  assign GEN_721 = {{2'd0}, 2'h2};
  assign T_7212 = T_7158_bpmatch & GEN_721;
  assign GEN_25 = T_7212;
  assign GEN_300 = 1'h0 == reg_tdrselect_tdrindex ? GEN_25 : GEN_284;
  assign GEN_327 = T_6267 ? GEN_300 : reg_bp_0_control_bpmatch;
  assign GEN_330 = T_6267 ? GEN_286 : reg_bp_0_control_m;
  assign GEN_336 = T_6267 ? GEN_290 : reg_bp_0_control_s;
  assign GEN_339 = T_6267 ? GEN_292 : reg_bp_0_control_u;
  assign GEN_342 = T_6267 ? GEN_294 : reg_bp_0_control_r;
  assign GEN_345 = T_6267 ? GEN_296 : reg_bp_0_control_w;
  assign GEN_348 = T_6267 ? GEN_298 : reg_bp_0_control_x;
  assign GEN_26 = wdata[38:0];
  assign GEN_351 = 1'h0 == reg_tdrselect_tdrindex ? GEN_26 : reg_bp_0_address;
  assign GEN_354 = T_6269 ? GEN_351 : reg_bp_0_address;
  assign GEN_381 = T_7131 ? GEN_327 : reg_bp_0_control_bpmatch;
  assign GEN_384 = T_7131 ? GEN_330 : reg_bp_0_control_m;
  assign GEN_390 = T_7131 ? GEN_336 : reg_bp_0_control_s;
  assign GEN_393 = T_7131 ? GEN_339 : reg_bp_0_control_u;
  assign GEN_396 = T_7131 ? GEN_342 : reg_bp_0_control_r;
  assign GEN_399 = T_7131 ? GEN_345 : reg_bp_0_control_w;
  assign GEN_402 = T_7131 ? GEN_348 : reg_bp_0_control_x;
  assign GEN_406 = T_7131 ? GEN_354 : reg_bp_0_address;
  assign GEN_432 = wen ? GEN_167 : GEN_135;
  assign GEN_433 = wen ? GEN_168 : GEN_136;
  assign GEN_434 = wen ? GEN_169 : reg_mstatus_mprv;
  assign GEN_435 = wen ? GEN_170 : GEN_137;
  assign GEN_436 = wen ? GEN_250 : reg_mstatus_pum;
  assign GEN_437 = wen ? GEN_249 : GEN_132;
  assign GEN_438 = wen ? GEN_248 : GEN_131;
  assign GEN_439 = wen ? GEN_247 : GEN_130;
  assign GEN_440 = wen ? GEN_175 : reg_mstatus_vm;
  assign GEN_441 = wen ? GEN_251 : reg_mstatus_fs;
  assign GEN_455 = wen ? GEN_265 : reg_mip_ssip;
  assign GEN_456 = wen ? GEN_191 : reg_mip_stip;
  assign GEN_457 = wen ? GEN_266 : reg_mie;
  assign GEN_458 = wen ? GEN_193 : {{24'd0}, GEN_110};
  assign GEN_459 = wen ? GEN_194 : reg_mscratch;
  assign GEN_460 = wen ? GEN_195 : {{32'd0}, reg_mtvec};
  assign GEN_461 = wen ? GEN_196 : GEN_111;
  assign GEN_462 = wen ? GEN_197 : GEN_112;
  assign GEN_480 = wen ? GEN_215 : reg_dcsr_halt;
  assign GEN_481 = wen ? GEN_216 : reg_dcsr_step;
  assign GEN_482 = wen ? GEN_217 : reg_dcsr_ebreakm;
  assign GEN_483 = wen ? GEN_218 : reg_dcsr_ebreaks;
  assign GEN_484 = wen ? GEN_219 : reg_dcsr_ebreaku;
  assign GEN_485 = wen ? GEN_220 : GEN_102;
  assign GEN_486 = wen ? GEN_221 : {{24'd0}, GEN_100};
  assign GEN_487 = wen ? GEN_222 : reg_dscratch;
  assign GEN_525 = wen ? GEN_267 : reg_sscratch;
  assign GEN_526 = wen ? GEN_268 : reg_sptbr_ppn;
  assign GEN_527 = wen ? GEN_269 : {{24'd0}, GEN_103};
  assign GEN_528 = wen ? GEN_270 : {{25'd0}, reg_stvec};
  assign GEN_529 = wen ? GEN_271 : GEN_104;
  assign GEN_530 = wen ? GEN_272 : GEN_105;
  assign GEN_531 = wen ? GEN_273 : reg_mideleg;
  assign GEN_532 = wen ? GEN_274 : reg_medeleg;
  assign GEN_536 = wen ? GEN_275 : reg_tdrselect_tdrindex;
  assign GEN_562 = wen ? GEN_381 : reg_bp_0_control_bpmatch;
  assign GEN_565 = wen ? GEN_384 : reg_bp_0_control_m;
  assign GEN_571 = wen ? GEN_390 : reg_bp_0_control_s;
  assign GEN_574 = wen ? GEN_393 : reg_bp_0_control_u;
  assign GEN_577 = wen ? GEN_396 : reg_bp_0_control_r;
  assign GEN_580 = wen ? GEN_399 : reg_bp_0_control_w;
  assign GEN_583 = wen ? GEN_402 : reg_bp_0_control_x;
  assign GEN_587 = wen ? GEN_406 : reg_bp_0_address;
  assign GEN_589 = reset ? 1'h0 : GEN_577;
  assign GEN_590 = reset ? 1'h0 : GEN_580;
  assign GEN_591 = reset ? 1'h0 : GEN_583;
  assign T_7278_control_tdrtype = T_7307;
  assign T_7278_control_bpamaskmax = T_7306;
  assign T_7278_control_reserved = T_7305;
  assign T_7278_control_bpaction = T_7304;
  assign T_7278_control_bpmatch = T_7303;
  assign T_7278_control_m = T_7302;
  assign T_7278_control_h = T_7301;
  assign T_7278_control_s = T_7300;
  assign T_7278_control_u = T_7299;
  assign T_7278_control_r = T_7298;
  assign T_7278_control_w = T_7297;
  assign T_7278_control_x = T_7296;
  assign T_7278_address = T_7295;
  assign T_7294 = {{102'd0}, 1'h0};
  assign T_7295 = T_7294[38:0];
  assign T_7296 = T_7294[39];
  assign T_7297 = T_7294[40];
  assign T_7298 = T_7294[41];
  assign T_7299 = T_7294[42];
  assign T_7300 = T_7294[43];
  assign T_7301 = T_7294[44];
  assign T_7302 = T_7294[45];
  assign T_7303 = T_7294[49:46];
  assign T_7304 = T_7294[57:50];
  assign T_7305 = T_7294[93:58];
  assign T_7306 = T_7294[98:94];
  assign T_7307 = T_7294[102:99];
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_235 = {1{$random}};
  reg_mstatus_debug = GEN_235[0:0];
  GEN_236 = {1{$random}};
  reg_mstatus_prv = GEN_236[1:0];
  GEN_237 = {1{$random}};
  reg_mstatus_sd = GEN_237[0:0];
  GEN_238 = {1{$random}};
  reg_mstatus_zero3 = GEN_238[30:0];
  GEN_239 = {1{$random}};
  reg_mstatus_sd_rv32 = GEN_239[0:0];
  GEN_240 = {1{$random}};
  reg_mstatus_zero2 = GEN_240[1:0];
  GEN_241 = {1{$random}};
  reg_mstatus_vm = GEN_241[4:0];
  GEN_242 = {1{$random}};
  reg_mstatus_zero1 = GEN_242[4:0];
  GEN_243 = {1{$random}};
  reg_mstatus_pum = GEN_243[0:0];
  GEN_244 = {1{$random}};
  reg_mstatus_mprv = GEN_244[0:0];
  GEN_245 = {1{$random}};
  reg_mstatus_xs = GEN_245[1:0];
  GEN_246 = {1{$random}};
  reg_mstatus_fs = GEN_246[1:0];
  GEN_252 = {1{$random}};
  reg_mstatus_mpp = GEN_252[1:0];
  GEN_253 = {1{$random}};
  reg_mstatus_hpp = GEN_253[1:0];
  GEN_254 = {1{$random}};
  reg_mstatus_spp = GEN_254[0:0];
  GEN_255 = {1{$random}};
  reg_mstatus_mpie = GEN_255[0:0];
  GEN_256 = {1{$random}};
  reg_mstatus_hpie = GEN_256[0:0];
  GEN_257 = {1{$random}};
  reg_mstatus_spie = GEN_257[0:0];
  GEN_258 = {1{$random}};
  reg_mstatus_upie = GEN_258[0:0];
  GEN_259 = {1{$random}};
  reg_mstatus_mie = GEN_259[0:0];
  GEN_260 = {1{$random}};
  reg_mstatus_hie = GEN_260[0:0];
  GEN_261 = {1{$random}};
  reg_mstatus_sie = GEN_261[0:0];
  GEN_262 = {1{$random}};
  reg_mstatus_uie = GEN_262[0:0];
  GEN_263 = {1{$random}};
  reg_dcsr_xdebugver = GEN_263[1:0];
  GEN_264 = {1{$random}};
  reg_dcsr_ndreset = GEN_264[0:0];
  GEN_276 = {1{$random}};
  reg_dcsr_fullreset = GEN_276[0:0];
  GEN_277 = {1{$random}};
  reg_dcsr_hwbpcount = GEN_277[11:0];
  GEN_278 = {1{$random}};
  reg_dcsr_ebreakm = GEN_278[0:0];
  GEN_279 = {1{$random}};
  reg_dcsr_ebreakh = GEN_279[0:0];
  GEN_280 = {1{$random}};
  reg_dcsr_ebreaks = GEN_280[0:0];
  GEN_281 = {1{$random}};
  reg_dcsr_ebreaku = GEN_281[0:0];
  GEN_282 = {1{$random}};
  reg_dcsr_zero2 = GEN_282[0:0];
  GEN_283 = {1{$random}};
  reg_dcsr_stopcycle = GEN_283[0:0];
  GEN_285 = {1{$random}};
  reg_dcsr_stoptime = GEN_285[0:0];
  GEN_287 = {1{$random}};
  reg_dcsr_cause = GEN_287[2:0];
  GEN_288 = {1{$random}};
  reg_dcsr_debugint = GEN_288[0:0];
  GEN_289 = {1{$random}};
  reg_dcsr_zero1 = GEN_289[0:0];
  GEN_291 = {1{$random}};
  reg_dcsr_halt = GEN_291[0:0];
  GEN_293 = {1{$random}};
  reg_dcsr_step = GEN_293[0:0];
  GEN_295 = {1{$random}};
  reg_dcsr_prv = GEN_295[1:0];
  GEN_297 = {1{$random}};
  reg_debug = GEN_297[0:0];
  GEN_299 = {2{$random}};
  reg_dpc = GEN_299[39:0];
  GEN_301 = {2{$random}};
  reg_dscratch = GEN_301[63:0];
  GEN_302 = {1{$random}};
  reg_singleStepped = GEN_302[0:0];
  GEN_303 = {1{$random}};
  reg_tdrselect_tdrmode = GEN_303[0:0];
  GEN_304 = {2{$random}};
  reg_tdrselect_reserved = GEN_304[61:0];
  GEN_305 = {1{$random}};
  reg_tdrselect_tdrindex = GEN_305[0:0];
  GEN_306 = {1{$random}};
  reg_bp_0_control_tdrtype = GEN_306[3:0];
  GEN_307 = {1{$random}};
  reg_bp_0_control_bpamaskmax = GEN_307[4:0];
  GEN_308 = {2{$random}};
  reg_bp_0_control_reserved = GEN_308[35:0];
  GEN_309 = {1{$random}};
  reg_bp_0_control_bpaction = GEN_309[7:0];
  GEN_310 = {1{$random}};
  reg_bp_0_control_bpmatch = GEN_310[3:0];
  GEN_311 = {1{$random}};
  reg_bp_0_control_m = GEN_311[0:0];
  GEN_312 = {1{$random}};
  reg_bp_0_control_h = GEN_312[0:0];
  GEN_313 = {1{$random}};
  reg_bp_0_control_s = GEN_313[0:0];
  GEN_314 = {1{$random}};
  reg_bp_0_control_u = GEN_314[0:0];
  GEN_315 = {1{$random}};
  reg_bp_0_control_r = GEN_315[0:0];
  GEN_316 = {1{$random}};
  reg_bp_0_control_w = GEN_316[0:0];
  GEN_317 = {1{$random}};
  reg_bp_0_control_x = GEN_317[0:0];
  GEN_318 = {2{$random}};
  reg_bp_0_address = GEN_318[38:0];
  GEN_319 = {1{$random}};
  reg_bp_1_control_tdrtype = GEN_319[3:0];
  GEN_320 = {1{$random}};
  reg_bp_1_control_bpamaskmax = GEN_320[4:0];
  GEN_321 = {2{$random}};
  reg_bp_1_control_reserved = GEN_321[35:0];
  GEN_322 = {1{$random}};
  reg_bp_1_control_bpaction = GEN_322[7:0];
  GEN_323 = {1{$random}};
  reg_bp_1_control_bpmatch = GEN_323[3:0];
  GEN_324 = {1{$random}};
  reg_bp_1_control_m = GEN_324[0:0];
  GEN_325 = {1{$random}};
  reg_bp_1_control_h = GEN_325[0:0];
  GEN_326 = {1{$random}};
  reg_bp_1_control_s = GEN_326[0:0];
  GEN_328 = {1{$random}};
  reg_bp_1_control_u = GEN_328[0:0];
  GEN_329 = {1{$random}};
  reg_bp_1_control_r = GEN_329[0:0];
  GEN_331 = {1{$random}};
  reg_bp_1_control_w = GEN_331[0:0];
  GEN_332 = {1{$random}};
  reg_bp_1_control_x = GEN_332[0:0];
  GEN_333 = {2{$random}};
  reg_bp_1_address = GEN_333[38:0];
  GEN_334 = {2{$random}};
  reg_mie = GEN_334[63:0];
  GEN_335 = {2{$random}};
  reg_mideleg = GEN_335[63:0];
  GEN_337 = {2{$random}};
  reg_medeleg = GEN_337[63:0];
  GEN_338 = {1{$random}};
  reg_mip_rocc = GEN_338[0:0];
  GEN_340 = {1{$random}};
  reg_mip_meip = GEN_340[0:0];
  GEN_341 = {1{$random}};
  reg_mip_heip = GEN_341[0:0];
  GEN_343 = {1{$random}};
  reg_mip_seip = GEN_343[0:0];
  GEN_344 = {1{$random}};
  reg_mip_ueip = GEN_344[0:0];
  GEN_346 = {1{$random}};
  reg_mip_mtip = GEN_346[0:0];
  GEN_347 = {1{$random}};
  reg_mip_htip = GEN_347[0:0];
  GEN_349 = {1{$random}};
  reg_mip_stip = GEN_349[0:0];
  GEN_350 = {1{$random}};
  reg_mip_utip = GEN_350[0:0];
  GEN_352 = {1{$random}};
  reg_mip_msip = GEN_352[0:0];
  GEN_353 = {1{$random}};
  reg_mip_hsip = GEN_353[0:0];
  GEN_355 = {1{$random}};
  reg_mip_ssip = GEN_355[0:0];
  GEN_356 = {1{$random}};
  reg_mip_usip = GEN_356[0:0];
  GEN_357 = {2{$random}};
  reg_mepc = GEN_357[39:0];
  GEN_358 = {2{$random}};
  reg_mcause = GEN_358[63:0];
  GEN_359 = {2{$random}};
  reg_mbadaddr = GEN_359[39:0];
  GEN_360 = {2{$random}};
  reg_mscratch = GEN_360[63:0];
  GEN_361 = {1{$random}};
  reg_mtvec = GEN_361[31:0];
  GEN_362 = {2{$random}};
  reg_sepc = GEN_362[39:0];
  GEN_363 = {2{$random}};
  reg_scause = GEN_363[63:0];
  GEN_364 = {2{$random}};
  reg_sbadaddr = GEN_364[39:0];
  GEN_365 = {2{$random}};
  reg_sscratch = GEN_365[63:0];
  GEN_366 = {2{$random}};
  reg_stvec = GEN_366[38:0];
  GEN_367 = {1{$random}};
  reg_sptbr_asid = GEN_367[6:0];
  GEN_368 = {2{$random}};
  reg_sptbr_ppn = GEN_368[37:0];
  GEN_369 = {1{$random}};
  reg_wfi = GEN_369[0:0];
  GEN_370 = {1{$random}};
  T_5544 = GEN_370[5:0];
  GEN_371 = {2{$random}};
  T_5552 = GEN_371[57:0];
  GEN_372 = {1{$random}};
  T_5560 = GEN_372[5:0];
  GEN_373 = {2{$random}};
  T_5568 = GEN_373[57:0];
  GEN_374 = {1{$random}};
  T_5576 = GEN_374[5:0];
  GEN_375 = {2{$random}};
  T_5584 = GEN_375[57:0];
  GEN_376 = {1{$random}};
  T_5592 = GEN_376[5:0];
  GEN_377 = {2{$random}};
  T_5600 = GEN_377[57:0];
  GEN_378 = {1{$random}};
  T_5608 = GEN_378[5:0];
  GEN_379 = {2{$random}};
  T_5616 = GEN_379[57:0];
  GEN_380 = {1{$random}};
  T_5624 = GEN_380[5:0];
  GEN_382 = {2{$random}};
  T_5632 = GEN_382[57:0];
  GEN_383 = {1{$random}};
  T_5640 = GEN_383[5:0];
  GEN_385 = {2{$random}};
  T_5648 = GEN_385[57:0];
  GEN_386 = {1{$random}};
  T_5656 = GEN_386[5:0];
  GEN_387 = {2{$random}};
  T_5664 = GEN_387[57:0];
  GEN_388 = {1{$random}};
  T_5672 = GEN_388[5:0];
  GEN_389 = {2{$random}};
  T_5680 = GEN_389[57:0];
  GEN_391 = {1{$random}};
  T_5688 = GEN_391[5:0];
  GEN_392 = {2{$random}};
  T_5696 = GEN_392[57:0];
  GEN_394 = {1{$random}};
  T_5704 = GEN_394[5:0];
  GEN_395 = {2{$random}};
  T_5712 = GEN_395[57:0];
  GEN_397 = {1{$random}};
  T_5720 = GEN_397[5:0];
  GEN_398 = {2{$random}};
  T_5728 = GEN_398[57:0];
  GEN_400 = {1{$random}};
  T_5736 = GEN_400[5:0];
  GEN_401 = {2{$random}};
  T_5744 = GEN_401[57:0];
  GEN_403 = {1{$random}};
  T_5752 = GEN_403[5:0];
  GEN_404 = {2{$random}};
  T_5760 = GEN_404[57:0];
  GEN_405 = {1{$random}};
  T_5768 = GEN_405[5:0];
  GEN_407 = {2{$random}};
  T_5776 = GEN_407[57:0];
  GEN_408 = {1{$random}};
  T_5784 = GEN_408[5:0];
  GEN_409 = {2{$random}};
  T_5792 = GEN_409[57:0];
  GEN_410 = {1{$random}};
  reg_fflags = GEN_410[4:0];
  GEN_411 = {1{$random}};
  reg_frm = GEN_411[2:0];
  GEN_412 = {1{$random}};
  T_5802 = GEN_412[5:0];
  GEN_413 = {2{$random}};
  T_5810 = GEN_413[57:0];
  GEN_414 = {1{$random}};
  T_5819 = GEN_414[5:0];
  GEN_415 = {2{$random}};
  T_5827 = GEN_415[57:0];
  GEN_416 = {1{$random}};
  GEN_63 = GEN_416[0:0];
  GEN_417 = {1{$random}};
  GEN_143 = GEN_417[6:0];
  GEN_418 = {1{$random}};
  GEN_144 = GEN_418[4:0];
  GEN_419 = {1{$random}};
  GEN_145 = GEN_419[4:0];
  GEN_420 = {1{$random}};
  GEN_146 = GEN_420[0:0];
  GEN_421 = {1{$random}};
  GEN_147 = GEN_421[0:0];
  GEN_422 = {1{$random}};
  GEN_148 = GEN_422[0:0];
  GEN_423 = {1{$random}};
  GEN_149 = GEN_423[4:0];
  GEN_424 = {1{$random}};
  GEN_150 = GEN_424[6:0];
  GEN_425 = {2{$random}};
  GEN_151 = GEN_425[63:0];
  GEN_426 = {2{$random}};
  GEN_152 = GEN_426[63:0];
  GEN_427 = {1{$random}};
  GEN_153 = GEN_427[0:0];
  GEN_428 = {1{$random}};
  GEN_154 = GEN_428[0:0];
  GEN_429 = {1{$random}};
  GEN_155 = GEN_429[0:0];
  GEN_430 = {1{$random}};
  GEN_156 = GEN_430[0:0];
  GEN_431 = {2{$random}};
  GEN_157 = GEN_431[39:0];
  GEN_442 = {1{$random}};
  GEN_158 = GEN_442[8:0];
  GEN_443 = {1{$random}};
  GEN_159 = GEN_443[4:0];
  GEN_444 = {1{$random}};
  GEN_160 = GEN_444[2:0];
  GEN_445 = {2{$random}};
  GEN_161 = GEN_445[63:0];
  GEN_446 = {1{$random}};
  GEN_162 = GEN_446[0:0];
  GEN_447 = {1{$random}};
  GEN_163 = GEN_447[0:0];
  GEN_448 = {2{$random}};
  GEN_164 = GEN_448[63:0];
  GEN_449 = {2{$random}};
  GEN_165 = GEN_449[63:0];
  GEN_450 = {1{$random}};
  GEN_166 = GEN_450[0:0];
  GEN_451 = {1{$random}};
  GEN_177 = GEN_451[0:0];
  GEN_452 = {1{$random}};
  GEN_178 = GEN_452[0:0];
  GEN_453 = {1{$random}};
  GEN_179 = GEN_453[0:0];
  GEN_454 = {1{$random}};
  GEN_180 = GEN_454[0:0];
  GEN_463 = {1{$random}};
  GEN_181 = GEN_463[0:0];
  GEN_464 = {1{$random}};
  GEN_182 = GEN_464[0:0];
  GEN_465 = {1{$random}};
  GEN_183 = GEN_465[1:0];
  GEN_466 = {1{$random}};
  GEN_184 = GEN_466[0:0];
  GEN_467 = {1{$random}};
  GEN_185 = GEN_467[30:0];
  GEN_468 = {1{$random}};
  GEN_186 = GEN_468[0:0];
  GEN_469 = {1{$random}};
  GEN_187 = GEN_469[1:0];
  GEN_470 = {1{$random}};
  GEN_188 = GEN_470[4:0];
  GEN_471 = {1{$random}};
  GEN_189 = GEN_471[4:0];
  GEN_472 = {1{$random}};
  GEN_198 = GEN_472[0:0];
  GEN_473 = {1{$random}};
  GEN_199 = GEN_473[0:0];
  GEN_474 = {1{$random}};
  GEN_200 = GEN_474[1:0];
  GEN_475 = {1{$random}};
  GEN_201 = GEN_475[1:0];
  GEN_476 = {1{$random}};
  GEN_202 = GEN_476[1:0];
  GEN_477 = {1{$random}};
  GEN_203 = GEN_477[1:0];
  GEN_478 = {1{$random}};
  GEN_204 = GEN_478[0:0];
  GEN_479 = {1{$random}};
  GEN_205 = GEN_479[0:0];
  GEN_488 = {1{$random}};
  GEN_206 = GEN_488[0:0];
  GEN_489 = {1{$random}};
  GEN_207 = GEN_489[0:0];
  GEN_490 = {1{$random}};
  GEN_208 = GEN_490[0:0];
  GEN_491 = {1{$random}};
  GEN_209 = GEN_491[0:0];
  GEN_492 = {1{$random}};
  GEN_210 = GEN_492[0:0];
  GEN_493 = {1{$random}};
  GEN_211 = GEN_493[0:0];
  GEN_494 = {1{$random}};
  GEN_212 = GEN_494[0:0];
  GEN_495 = {1{$random}};
  GEN_213 = GEN_495[0:0];
  GEN_496 = {1{$random}};
  GEN_214 = GEN_496[0:0];
  GEN_497 = {1{$random}};
  GEN_223 = GEN_497[2:0];
  GEN_498 = {1{$random}};
  GEN_224 = GEN_498[1:0];
  GEN_499 = {1{$random}};
  GEN_225 = GEN_499[2:0];
  GEN_500 = {1{$random}};
  GEN_226 = GEN_500[0:0];
  GEN_501 = {1{$random}};
  GEN_227 = GEN_501[3:0];
  GEN_502 = {2{$random}};
  GEN_228 = GEN_502[63:0];
  GEN_503 = {1{$random}};
  GEN_229 = GEN_503[0:0];
  GEN_504 = {1{$random}};
  GEN_230 = GEN_504[0:0];
  GEN_505 = {3{$random}};
  GEN_231 = GEN_505[64:0];
  GEN_506 = {1{$random}};
  GEN_232 = GEN_506[4:0];
  GEN_507 = {1{$random}};
  GEN_233 = GEN_507[0:0];
  GEN_508 = {1{$random}};
  GEN_234 = GEN_508[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      reg_mstatus_debug <= reset_mstatus_debug;
    end
    if(reset) begin
      reg_mstatus_prv <= reset_mstatus_prv;
    end else begin
      if(insn_ret) begin
        if(T_6536) begin
          reg_mstatus_prv <= reg_mstatus_mpp;
        end else begin
          if(T_6530) begin
            reg_mstatus_prv <= reg_dcsr_prv;
          end else begin
            if(T_6482) begin
              reg_mstatus_prv <= {{1'd0}, reg_mstatus_spp};
            end else begin
              if(exception) begin
                if(T_6517) begin
                  reg_mstatus_prv <= 2'h3;
                end else begin
                  if(T_6510) begin
                    reg_mstatus_prv <= {{1'd0}, 1'h1};
                  end
                end
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6517) begin
            reg_mstatus_prv <= 2'h3;
          end else begin
            if(T_6510) begin
              reg_mstatus_prv <= {{1'd0}, 1'h1};
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_sd <= reset_mstatus_sd;
    end
    if(reset) begin
      reg_mstatus_zero3 <= reset_mstatus_zero3;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= reset_mstatus_sd_rv32;
    end
    if(reset) begin
      reg_mstatus_zero2 <= reset_mstatus_zero2;
    end
    if(reset) begin
      reg_mstatus_vm <= reset_mstatus_vm;
    end else begin
      if(wen) begin
        if(T_6291) begin
          if(T_6798) begin
            reg_mstatus_vm <= {{1'd0}, 4'h9};
          end else begin
            if(T_6795) begin
              reg_mstatus_vm <= {{4'd0}, 1'h0};
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_zero1 <= reset_mstatus_zero1;
    end
    if(reset) begin
      reg_mstatus_pum <= reset_mstatus_pum;
    end else begin
      if(wen) begin
        if(T_6319) begin
          reg_mstatus_pum <= T_6993_pum;
        end else begin
          if(T_6291) begin
            reg_mstatus_pum <= T_6738_pum;
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_mprv <= reset_mstatus_mprv;
    end else begin
      if(wen) begin
        if(T_6291) begin
          reg_mstatus_mprv <= T_6738_mprv;
        end
      end
    end
    if(reset) begin
      reg_mstatus_xs <= reset_mstatus_xs;
    end
    if(reset) begin
      reg_mstatus_fs <= reset_mstatus_fs;
    end else begin
      if(wen) begin
        if(T_6319) begin
          reg_mstatus_fs <= T_7046;
        end else begin
          if(T_6291) begin
            reg_mstatus_fs <= T_6804;
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_mpp <= reset_mstatus_mpp;
    end else begin
      if(wen) begin
        if(T_6291) begin
          if(T_6793) begin
            reg_mstatus_mpp <= T_6738_mpp;
          end else begin
            if(insn_ret) begin
              if(T_6536) begin
                reg_mstatus_mpp <= {{1'd0}, 1'h0};
              end else begin
                if(exception) begin
                  if(T_6517) begin
                    reg_mstatus_mpp <= reg_mstatus_prv;
                  end
                end
              end
            end else begin
              if(exception) begin
                if(T_6517) begin
                  reg_mstatus_mpp <= reg_mstatus_prv;
                end
              end
            end
          end
        end else begin
          if(insn_ret) begin
            if(T_6536) begin
              reg_mstatus_mpp <= {{1'd0}, 1'h0};
            end else begin
              if(exception) begin
                if(T_6517) begin
                  reg_mstatus_mpp <= reg_mstatus_prv;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6517) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6536) begin
            reg_mstatus_mpp <= {{1'd0}, 1'h0};
          end else begin
            reg_mstatus_mpp <= GEN_114;
          end
        end else begin
          reg_mstatus_mpp <= GEN_114;
        end
      end
    end
    if(reset) begin
      reg_mstatus_hpp <= reset_mstatus_hpp;
    end
    if(reset) begin
      reg_mstatus_spp <= reset_mstatus_spp;
    end else begin
      reg_mstatus_spp <= GEN_437[0];
    end
    if(reset) begin
      reg_mstatus_mpie <= reset_mstatus_mpie;
    end else begin
      if(wen) begin
        if(T_6291) begin
          reg_mstatus_mpie <= T_6738_mpie;
        end else begin
          if(insn_ret) begin
            if(T_6536) begin
              reg_mstatus_mpie <= 1'h0;
            end else begin
              if(exception) begin
                if(T_6517) begin
                  reg_mstatus_mpie <= T_6501;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6517) begin
                reg_mstatus_mpie <= T_6501;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6536) begin
            reg_mstatus_mpie <= 1'h0;
          end else begin
            if(exception) begin
              if(T_6517) begin
                reg_mstatus_mpie <= T_6501;
              end
            end
          end
        end else begin
          if(exception) begin
            if(T_6517) begin
              reg_mstatus_mpie <= T_6501;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_hpie <= reset_mstatus_hpie;
    end
    if(reset) begin
      reg_mstatus_spie <= reset_mstatus_spie;
    end else begin
      if(wen) begin
        if(T_6319) begin
          reg_mstatus_spie <= T_6993_spie;
        end else begin
          if(T_6291) begin
            reg_mstatus_spie <= T_6738_spie;
          end else begin
            if(insn_ret) begin
              if(T_6482) begin
                reg_mstatus_spie <= 1'h0;
              end else begin
                if(exception) begin
                  if(T_6510) begin
                    reg_mstatus_spie <= T_6501;
                  end
                end
              end
            end else begin
              if(exception) begin
                if(T_6510) begin
                  reg_mstatus_spie <= T_6501;
                end
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6482) begin
            reg_mstatus_spie <= 1'h0;
          end else begin
            if(exception) begin
              if(T_6510) begin
                reg_mstatus_spie <= T_6501;
              end
            end
          end
        end else begin
          if(exception) begin
            if(T_6510) begin
              reg_mstatus_spie <= T_6501;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_upie <= reset_mstatus_upie;
    end
    if(reset) begin
      reg_mstatus_mie <= reset_mstatus_mie;
    end else begin
      if(wen) begin
        if(T_6291) begin
          reg_mstatus_mie <= T_6738_mie;
        end else begin
          if(insn_ret) begin
            if(T_6536) begin
              if(T_6537) begin
                reg_mstatus_mie <= reg_mstatus_mpie;
              end else begin
                if(exception) begin
                  if(T_6517) begin
                    reg_mstatus_mie <= 1'h0;
                  end
                end
              end
            end else begin
              if(exception) begin
                if(T_6517) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6517) begin
                reg_mstatus_mie <= 1'h0;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6536) begin
            if(T_6537) begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end else begin
              if(exception) begin
                if(T_6517) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            reg_mstatus_mie <= GEN_115;
          end
        end else begin
          reg_mstatus_mie <= GEN_115;
        end
      end
    end
    if(reset) begin
      reg_mstatus_hie <= reset_mstatus_hie;
    end
    if(reset) begin
      reg_mstatus_sie <= reset_mstatus_sie;
    end else begin
      if(wen) begin
        if(T_6319) begin
          reg_mstatus_sie <= T_6993_sie;
        end else begin
          if(T_6291) begin
            reg_mstatus_sie <= T_6738_sie;
          end else begin
            if(insn_ret) begin
              if(T_6536) begin
                if(T_6543) begin
                  reg_mstatus_sie <= reg_mstatus_mpie;
                end else begin
                  if(T_6482) begin
                    if(reg_mstatus_spp) begin
                      reg_mstatus_sie <= reg_mstatus_spie;
                    end else begin
                      if(exception) begin
                        if(T_6510) begin
                          reg_mstatus_sie <= 1'h0;
                        end
                      end
                    end
                  end else begin
                    if(exception) begin
                      if(T_6510) begin
                        reg_mstatus_sie <= 1'h0;
                      end
                    end
                  end
                end
              end else begin
                if(T_6482) begin
                  if(reg_mstatus_spp) begin
                    reg_mstatus_sie <= reg_mstatus_spie;
                  end else begin
                    if(exception) begin
                      if(T_6510) begin
                        reg_mstatus_sie <= 1'h0;
                      end
                    end
                  end
                end else begin
                  if(exception) begin
                    if(T_6510) begin
                      reg_mstatus_sie <= 1'h0;
                    end
                  end
                end
              end
            end else begin
              reg_mstatus_sie <= GEN_108;
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6536) begin
            if(T_6543) begin
              reg_mstatus_sie <= reg_mstatus_mpie;
            end else begin
              if(T_6482) begin
                if(reg_mstatus_spp) begin
                  reg_mstatus_sie <= reg_mstatus_spie;
                end else begin
                  reg_mstatus_sie <= GEN_108;
                end
              end else begin
                reg_mstatus_sie <= GEN_108;
              end
            end
          end else begin
            if(T_6482) begin
              if(reg_mstatus_spp) begin
                reg_mstatus_sie <= reg_mstatus_spie;
              end else begin
                reg_mstatus_sie <= GEN_108;
              end
            end else begin
              reg_mstatus_sie <= GEN_108;
            end
          end
        end else begin
          reg_mstatus_sie <= GEN_108;
        end
      end
    end
    if(reset) begin
      reg_mstatus_uie <= reset_mstatus_uie;
    end
    if(reset) begin
      reg_dcsr_xdebugver <= reset_dcsr_xdebugver;
    end
    if(reset) begin
      reg_dcsr_ndreset <= reset_dcsr_ndreset;
    end
    if(reset) begin
      reg_dcsr_fullreset <= reset_dcsr_fullreset;
    end
    if(reset) begin
      reg_dcsr_hwbpcount <= reset_dcsr_hwbpcount;
    end else begin
      reg_dcsr_hwbpcount <= {{11'd0}, 1'h1};
    end
    if(reset) begin
      reg_dcsr_ebreakm <= reset_dcsr_ebreakm;
    end else begin
      if(wen) begin
        if(T_6313) begin
          reg_dcsr_ebreakm <= T_6906_ebreakm;
        end
      end
    end
    if(reset) begin
      reg_dcsr_ebreakh <= reset_dcsr_ebreakh;
    end
    if(reset) begin
      reg_dcsr_ebreaks <= reset_dcsr_ebreaks;
    end else begin
      if(wen) begin
        if(T_6313) begin
          reg_dcsr_ebreaks <= T_6906_ebreaks;
        end
      end
    end
    if(reset) begin
      reg_dcsr_ebreaku <= reset_dcsr_ebreaku;
    end else begin
      if(wen) begin
        if(T_6313) begin
          reg_dcsr_ebreaku <= T_6906_ebreaku;
        end
      end
    end
    if(reset) begin
      reg_dcsr_zero2 <= reset_dcsr_zero2;
    end
    if(reset) begin
      reg_dcsr_stopcycle <= reset_dcsr_stopcycle;
    end
    if(reset) begin
      reg_dcsr_stoptime <= reset_dcsr_stoptime;
    end
    if(reset) begin
      reg_dcsr_cause <= reset_dcsr_cause;
    end else begin
      if(exception) begin
        if(T_6463) begin
          if(reg_singleStepped) begin
            reg_dcsr_cause <= 3'h4;
          end else begin
            reg_dcsr_cause <= {{1'd0}, T_6506};
          end
        end
      end
    end
    if(reset) begin
      reg_dcsr_debugint <= reset_dcsr_debugint;
    end else begin
      reg_dcsr_debugint <= io_prci_interrupts_debug;
    end
    if(reset) begin
      reg_dcsr_zero1 <= reset_dcsr_zero1;
    end
    if(reset) begin
      reg_dcsr_halt <= reset_dcsr_halt;
    end else begin
      if(wen) begin
        if(T_6313) begin
          reg_dcsr_halt <= T_6906_halt;
        end
      end
    end
    if(reset) begin
      reg_dcsr_step <= reset_dcsr_step;
    end else begin
      if(wen) begin
        if(T_6313) begin
          reg_dcsr_step <= T_6906_step;
        end
      end
    end
    if(reset) begin
      reg_dcsr_prv <= reset_dcsr_prv;
    end else begin
      if(wen) begin
        if(T_6313) begin
          reg_dcsr_prv <= T_6906_prv;
        end else begin
          if(exception) begin
            if(T_6463) begin
              reg_dcsr_prv <= reg_mstatus_prv;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6463) begin
            reg_dcsr_prv <= reg_mstatus_prv;
          end
        end
      end
    end
    if(reset) begin
      reg_debug <= 1'h0;
    end else begin
      if(insn_ret) begin
        if(T_6530) begin
          reg_debug <= 1'h0;
        end else begin
          if(exception) begin
            if(T_6463) begin
              reg_debug <= 1'h1;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6463) begin
            reg_debug <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_dpc <= GEN_486[39:0];
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6317) begin
          reg_dscratch <= wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5325) begin
        reg_singleStepped <= 1'h0;
      end else begin
        if(T_5322) begin
          reg_singleStepped <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_tdrselect_tdrmode <= 1'h1;
    end
    if(1'h0) begin
    end else begin
      reg_tdrselect_reserved <= {{61'd0}, 1'h0};
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6265) begin
          reg_tdrselect_tdrindex <= T_7124_tdrindex;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_tdrtype <= {{3'd0}, 1'h1};
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_bpamaskmax <= {{2'd0}, 3'h4};
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_reserved <= {{35'd0}, 1'h0};
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_bpaction <= {{7'd0}, 1'h0};
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7131) begin
          if(T_6267) begin
            if(1'h0 == reg_tdrselect_tdrindex) begin
              reg_bp_0_control_bpmatch <= GEN_25;
            end else begin
              if(1'h0 == reg_tdrselect_tdrindex) begin
                reg_bp_0_control_bpmatch <= GEN_17;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7131) begin
          if(T_6267) begin
            if(1'h0 == reg_tdrselect_tdrindex) begin
              reg_bp_0_control_m <= GEN_18;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_h <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7131) begin
          if(T_6267) begin
            if(1'h0 == reg_tdrselect_tdrindex) begin
              reg_bp_0_control_s <= GEN_20;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7131) begin
          if(T_6267) begin
            if(1'h0 == reg_tdrselect_tdrindex) begin
              reg_bp_0_control_u <= GEN_21;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_r <= 1'h0;
      end else begin
        if(wen) begin
          if(T_7131) begin
            if(T_6267) begin
              if(1'h0 == reg_tdrselect_tdrindex) begin
                reg_bp_0_control_r <= GEN_22;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_w <= 1'h0;
      end else begin
        if(wen) begin
          if(T_7131) begin
            if(T_6267) begin
              if(1'h0 == reg_tdrselect_tdrindex) begin
                reg_bp_0_control_w <= GEN_23;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_x <= 1'h0;
      end else begin
        if(wen) begin
          if(T_7131) begin
            if(T_6267) begin
              if(1'h0 == reg_tdrselect_tdrindex) begin
                reg_bp_0_control_x <= GEN_24;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7131) begin
          if(T_6269) begin
            if(1'h0 == reg_tdrselect_tdrindex) begin
              reg_bp_0_address <= GEN_26;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_tdrtype <= T_7278_control_tdrtype;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_bpamaskmax <= T_7278_control_bpamaskmax;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_reserved <= T_7278_control_reserved;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_bpaction <= T_7278_control_bpaction;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_bpmatch <= T_7278_control_bpmatch;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_m <= T_7278_control_m;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_h <= T_7278_control_h;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_s <= T_7278_control_s;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_u <= T_7278_control_u;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_r <= T_7278_control_r;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_w <= T_7278_control_w;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_x <= T_7278_control_x;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_address <= T_7278_address;
    end
    if(reset) begin
      reg_mie <= 64'h0;
    end else begin
      if(wen) begin
        if(T_6323) begin
          reg_mie <= T_7105;
        end else begin
          if(T_6297) begin
            reg_mie <= T_6860;
          end
        end
      end
    end
    if(reset) begin
      reg_mideleg <= 64'h0;
    end else begin
      if(wen) begin
        if(T_6299) begin
          reg_mideleg <= T_7114;
        end
      end
    end
    if(reset) begin
      reg_medeleg <= 64'h0;
    end else begin
      if(wen) begin
        if(T_6301) begin
          reg_medeleg <= T_7115;
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_meip <= io_prci_interrupts_meip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_seip <= io_prci_interrupts_seip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_mtip <= io_prci_interrupts_mtip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6295) begin
          reg_mip_stip <= T_6833_stip;
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_msip <= io_prci_interrupts_msip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6321) begin
          reg_mip_ssip <= T_7075_ssip;
        end else begin
          if(T_6295) begin
            reg_mip_ssip <= T_6833_ssip;
          end
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mepc <= GEN_458[39:0];
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6309) begin
          reg_mcause <= T_6868;
        end else begin
          if(exception) begin
            if(T_6517) begin
              if(T_6442) begin
                reg_mcause <= io_cause;
              end else begin
                reg_mcause <= {{60'd0}, T_6449};
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6517) begin
            if(T_6442) begin
              reg_mcause <= io_cause;
            end else begin
              reg_mcause <= {{60'd0}, T_6449};
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6307) begin
          reg_mbadaddr <= T_6869;
        end else begin
          if(exception) begin
            if(T_6517) begin
              reg_mbadaddr <= io_badaddr;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6517) begin
            reg_mbadaddr <= io_badaddr;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6303) begin
          reg_mscratch <= wdata;
        end
      end
    end
    if(reset) begin
      reg_mtvec <= 32'h1010;
    end else begin
      reg_mtvec <= GEN_460[31:0];
    end
    if(1'h0) begin
    end else begin
      reg_sepc <= GEN_527[39:0];
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6327) begin
          reg_scause <= T_6868;
        end else begin
          if(exception) begin
            if(T_6510) begin
              if(T_6442) begin
                reg_scause <= io_cause;
              end else begin
                reg_scause <= {{60'd0}, T_6449};
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6510) begin
            if(T_6442) begin
              reg_scause <= io_cause;
            end else begin
              reg_scause <= {{60'd0}, T_6449};
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6329) begin
          reg_sbadaddr <= T_6869;
        end else begin
          if(exception) begin
            if(T_6510) begin
              reg_sbadaddr <= io_badaddr;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6510) begin
            reg_sbadaddr <= io_badaddr;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6325) begin
          reg_sscratch <= wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_stvec <= GEN_528[38:0];
    end
    if(1'h0) begin
    end else begin
      reg_sptbr_asid <= {{6'd0}, 1'h0};
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6331) begin
          reg_sptbr_ppn <= {{18'd0}, T_7106};
        end
      end
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else begin
      if(T_6439) begin
        reg_wfi <= 1'h0;
      end else begin
        if(insn_wfi) begin
          reg_wfi <= 1'h1;
        end
      end
    end
    if(reset) begin
      T_5544 <= 6'h0;
    end else begin
      if(io_uarch_counters_0) begin
        T_5544 <= T_5550;
      end
    end
    if(reset) begin
      T_5552 <= 58'h0;
    end else begin
      if(T_5554) begin
        T_5552 <= T_5557;
      end
    end
    if(reset) begin
      T_5560 <= 6'h0;
    end else begin
      if(io_uarch_counters_1) begin
        T_5560 <= T_5566;
      end
    end
    if(reset) begin
      T_5568 <= 58'h0;
    end else begin
      if(T_5570) begin
        T_5568 <= T_5573;
      end
    end
    if(reset) begin
      T_5576 <= 6'h0;
    end else begin
      if(io_uarch_counters_2) begin
        T_5576 <= T_5582;
      end
    end
    if(reset) begin
      T_5584 <= 58'h0;
    end else begin
      if(T_5586) begin
        T_5584 <= T_5589;
      end
    end
    if(reset) begin
      T_5592 <= 6'h0;
    end else begin
      if(io_uarch_counters_3) begin
        T_5592 <= T_5598;
      end
    end
    if(reset) begin
      T_5600 <= 58'h0;
    end else begin
      if(T_5602) begin
        T_5600 <= T_5605;
      end
    end
    if(reset) begin
      T_5608 <= 6'h0;
    end else begin
      if(io_uarch_counters_4) begin
        T_5608 <= T_5614;
      end
    end
    if(reset) begin
      T_5616 <= 58'h0;
    end else begin
      if(T_5618) begin
        T_5616 <= T_5621;
      end
    end
    if(reset) begin
      T_5624 <= 6'h0;
    end else begin
      if(io_uarch_counters_5) begin
        T_5624 <= T_5630;
      end
    end
    if(reset) begin
      T_5632 <= 58'h0;
    end else begin
      if(T_5634) begin
        T_5632 <= T_5637;
      end
    end
    if(reset) begin
      T_5640 <= 6'h0;
    end else begin
      if(io_uarch_counters_6) begin
        T_5640 <= T_5646;
      end
    end
    if(reset) begin
      T_5648 <= 58'h0;
    end else begin
      if(T_5650) begin
        T_5648 <= T_5653;
      end
    end
    if(reset) begin
      T_5656 <= 6'h0;
    end else begin
      if(io_uarch_counters_7) begin
        T_5656 <= T_5662;
      end
    end
    if(reset) begin
      T_5664 <= 58'h0;
    end else begin
      if(T_5666) begin
        T_5664 <= T_5669;
      end
    end
    if(reset) begin
      T_5672 <= 6'h0;
    end else begin
      if(io_uarch_counters_8) begin
        T_5672 <= T_5678;
      end
    end
    if(reset) begin
      T_5680 <= 58'h0;
    end else begin
      if(T_5682) begin
        T_5680 <= T_5685;
      end
    end
    if(reset) begin
      T_5688 <= 6'h0;
    end else begin
      if(io_uarch_counters_9) begin
        T_5688 <= T_5694;
      end
    end
    if(reset) begin
      T_5696 <= 58'h0;
    end else begin
      if(T_5698) begin
        T_5696 <= T_5701;
      end
    end
    if(reset) begin
      T_5704 <= 6'h0;
    end else begin
      if(io_uarch_counters_10) begin
        T_5704 <= T_5710;
      end
    end
    if(reset) begin
      T_5712 <= 58'h0;
    end else begin
      if(T_5714) begin
        T_5712 <= T_5717;
      end
    end
    if(reset) begin
      T_5720 <= 6'h0;
    end else begin
      if(io_uarch_counters_11) begin
        T_5720 <= T_5726;
      end
    end
    if(reset) begin
      T_5728 <= 58'h0;
    end else begin
      if(T_5730) begin
        T_5728 <= T_5733;
      end
    end
    if(reset) begin
      T_5736 <= 6'h0;
    end else begin
      if(io_uarch_counters_12) begin
        T_5736 <= T_5742;
      end
    end
    if(reset) begin
      T_5744 <= 58'h0;
    end else begin
      if(T_5746) begin
        T_5744 <= T_5749;
      end
    end
    if(reset) begin
      T_5752 <= 6'h0;
    end else begin
      if(io_uarch_counters_13) begin
        T_5752 <= T_5758;
      end
    end
    if(reset) begin
      T_5760 <= 58'h0;
    end else begin
      if(T_5762) begin
        T_5760 <= T_5765;
      end
    end
    if(reset) begin
      T_5768 <= 6'h0;
    end else begin
      if(io_uarch_counters_14) begin
        T_5768 <= T_5774;
      end
    end
    if(reset) begin
      T_5776 <= 58'h0;
    end else begin
      if(T_5778) begin
        T_5776 <= T_5781;
      end
    end
    if(reset) begin
      T_5784 <= 6'h0;
    end else begin
      if(io_uarch_counters_15) begin
        T_5784 <= T_5790;
      end
    end
    if(reset) begin
      T_5792 <= 58'h0;
    end else begin
      if(T_5794) begin
        T_5792 <= T_5797;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_fcsr_flags_valid) begin
        reg_fflags <= T_6680;
      end
    end
    if(1'h0) begin
    end
    if(reset) begin
      T_5802 <= 6'h0;
    end else begin
      if(io_retire) begin
        T_5802 <= T_5808;
      end
    end
    if(reset) begin
      T_5810 <= 58'h0;
    end else begin
      if(T_5812) begin
        T_5810 <= T_5815;
      end
    end
    if(reset) begin
      T_5819 <= 6'h0;
    end else begin
      T_5819 <= T_5825;
    end
    if(reset) begin
      T_5827 <= 58'h0;
    end else begin
      if(T_5828) begin
        T_5827 <= T_5832;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at csr.scala:185 assert(!io.singleStep || io.retire <= UInt(1))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_5342) begin
          $fwrite(32'h80000002,"Assertion failed\n    at csr.scala:186 assert(!reg_singleStepped || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_5342) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_5342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_6558) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at csr.scala:442 assert(PopCount(insn_ret :: io.exception :: io.csr_xcpt :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_6558) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_6558) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BreakpointUnit(
  input   clk,
  input   reset,
  input   io_status_debug,
  input  [1:0] io_status_prv,
  input   io_status_sd,
  input  [30:0] io_status_zero3,
  input   io_status_sd_rv32,
  input  [1:0] io_status_zero2,
  input  [4:0] io_status_vm,
  input  [4:0] io_status_zero1,
  input   io_status_pum,
  input   io_status_mprv,
  input  [1:0] io_status_xs,
  input  [1:0] io_status_fs,
  input  [1:0] io_status_mpp,
  input  [1:0] io_status_hpp,
  input   io_status_spp,
  input   io_status_mpie,
  input   io_status_hpie,
  input   io_status_spie,
  input   io_status_upie,
  input   io_status_mie,
  input   io_status_hie,
  input   io_status_sie,
  input   io_status_uie,
  input  [3:0] io_bp_0_control_tdrtype,
  input  [4:0] io_bp_0_control_bpamaskmax,
  input  [35:0] io_bp_0_control_reserved,
  input  [7:0] io_bp_0_control_bpaction,
  input  [3:0] io_bp_0_control_bpmatch,
  input   io_bp_0_control_m,
  input   io_bp_0_control_h,
  input   io_bp_0_control_s,
  input   io_bp_0_control_u,
  input   io_bp_0_control_r,
  input   io_bp_0_control_w,
  input   io_bp_0_control_x,
  input  [38:0] io_bp_0_address,
  input  [38:0] io_pc,
  input  [38:0] io_ea,
  output  io_xcpt_if,
  output  io_xcpt_ld,
  output  io_xcpt_st
);
  wire [1:0] T_176;
  wire [1:0] T_177;
  wire [3:0] T_178;
  wire [3:0] T_179;
  wire  T_180;
  wire [38:0] T_181;
  wire  T_182;
  wire  T_184;
  wire  T_185;
  wire [1:0] T_186;
  wire  T_187;
  wire  T_188;
  wire  T_189;
  wire [2:0] T_190;
  wire  T_191;
  wire  T_192;
  wire  T_193;
  wire [3:0] T_194;
  wire [38:0] GEN_6;
  wire [38:0] T_195;
  wire [38:0] T_196;
  wire [38:0] T_210;
  wire  T_211;
  wire  T_212;
  wire [38:0] T_214;
  wire [38:0] T_228;
  wire  T_244;
  wire  T_245;
  wire  T_278;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  assign io_xcpt_if = GEN_3;
  assign io_xcpt_ld = GEN_4;
  assign io_xcpt_st = GEN_5;
  assign T_176 = {io_bp_0_control_s,io_bp_0_control_u};
  assign T_177 = {io_bp_0_control_m,io_bp_0_control_h};
  assign T_178 = {T_177,T_176};
  assign T_179 = T_178 >> io_status_prv;
  assign T_180 = T_179[0];
  assign T_181 = ~ io_pc;
  assign T_182 = io_bp_0_control_bpmatch[1];
  assign T_184 = io_bp_0_address[0];
  assign T_185 = T_182 & T_184;
  assign T_186 = {T_185,T_182};
  assign T_187 = T_186[1];
  assign T_188 = io_bp_0_address[1];
  assign T_189 = T_187 & T_188;
  assign T_190 = {T_189,T_186};
  assign T_191 = T_190[2];
  assign T_192 = io_bp_0_address[2];
  assign T_193 = T_191 & T_192;
  assign T_194 = {T_193,T_190};
  assign GEN_6 = {{35'd0}, T_194};
  assign T_195 = T_181 | GEN_6;
  assign T_196 = ~ io_bp_0_address;
  assign T_210 = T_196 | GEN_6;
  assign T_211 = T_195 == T_210;
  assign T_212 = T_211 & io_bp_0_control_x;
  assign T_214 = ~ io_ea;
  assign T_228 = T_214 | GEN_6;
  assign T_244 = T_228 == T_210;
  assign T_245 = T_244 & io_bp_0_control_r;
  assign T_278 = T_244 & io_bp_0_control_w;
  assign GEN_3 = T_180 ? T_212 : 1'h0;
  assign GEN_4 = T_180 ? T_245 : 1'h0;
  assign GEN_5 = T_180 ? T_278 : 1'h0;
endmodule
module ALU(
  input   clk,
  input   reset,
  input   io_dw,
  input  [3:0] io_fn,
  input  [63:0] io_in2,
  input  [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output  io_cmp_out
);
  wire  T_7;
  wire [63:0] T_8;
  wire [63:0] in2_inv;
  wire [63:0] in1_xor_in2;
  wire [64:0] T_9;
  wire [63:0] T_10;
  wire [63:0] GEN_1;
  wire [64:0] T_12;
  wire [63:0] T_13;
  wire  T_14;
  wire  T_17;
  wire [63:0] GEN_2;
  wire  T_19;
  wire  T_20;
  wire  T_21;
  wire  T_22;
  wire  T_23;
  wire  T_24;
  wire  T_27;
  wire  T_28;
  wire  T_29;
  wire  T_30;
  wire  T_32;
  wire  T_33;
  wire [31:0] GEN_3;
  wire [32:0] T_35;
  wire [31:0] T_36;
  wire [31:0] T_41;
  wire [31:0] T_42;
  wire  T_43;
  wire  T_48;
  wire [4:0] T_49;
  wire [5:0] shamt;
  wire [31:0] T_50;
  wire [63:0] shin_r;
  wire [3:0] GEN_4;
  wire  T_51;
  wire  T_52;
  wire  T_53;
  wire [31:0] T_58;
  wire [63:0] GEN_5;
  wire [63:0] T_59;
  wire [31:0] T_60;
  wire [63:0] GEN_6;
  wire [63:0] T_61;
  wire [63:0] T_63;
  wire [63:0] T_64;
  wire [47:0] T_68;
  wire [63:0] GEN_7;
  wire [63:0] T_69;
  wire [47:0] T_70;
  wire [63:0] GEN_8;
  wire [63:0] T_71;
  wire [63:0] T_73;
  wire [63:0] T_74;
  wire [55:0] T_78;
  wire [63:0] GEN_9;
  wire [63:0] T_79;
  wire [55:0] T_80;
  wire [63:0] GEN_10;
  wire [63:0] T_81;
  wire [63:0] T_83;
  wire [63:0] T_84;
  wire [59:0] T_88;
  wire [63:0] GEN_11;
  wire [63:0] T_89;
  wire [59:0] T_90;
  wire [63:0] GEN_12;
  wire [63:0] T_91;
  wire [63:0] T_93;
  wire [63:0] T_94;
  wire [61:0] T_98;
  wire [63:0] GEN_13;
  wire [63:0] T_99;
  wire [61:0] T_100;
  wire [63:0] GEN_14;
  wire [63:0] T_101;
  wire [63:0] T_103;
  wire [63:0] T_104;
  wire [62:0] T_108;
  wire [63:0] GEN_15;
  wire [63:0] T_109;
  wire [62:0] T_110;
  wire [63:0] GEN_16;
  wire [63:0] T_111;
  wire [63:0] T_113;
  wire [63:0] T_114;
  wire [63:0] shin;
  wire  T_116;
  wire  T_117;
  wire [64:0] T_118;
  wire [64:0] T_119;
  wire [64:0] T_120;
  wire [63:0] shout_r;
  wire [31:0] T_125;
  wire [63:0] GEN_17;
  wire [63:0] T_126;
  wire [31:0] T_127;
  wire [63:0] GEN_18;
  wire [63:0] T_128;
  wire [63:0] T_130;
  wire [63:0] T_131;
  wire [47:0] T_135;
  wire [63:0] GEN_19;
  wire [63:0] T_136;
  wire [47:0] T_137;
  wire [63:0] GEN_20;
  wire [63:0] T_138;
  wire [63:0] T_140;
  wire [63:0] T_141;
  wire [55:0] T_145;
  wire [63:0] GEN_21;
  wire [63:0] T_146;
  wire [55:0] T_147;
  wire [63:0] GEN_22;
  wire [63:0] T_148;
  wire [63:0] T_150;
  wire [63:0] T_151;
  wire [59:0] T_155;
  wire [63:0] GEN_23;
  wire [63:0] T_156;
  wire [59:0] T_157;
  wire [63:0] GEN_24;
  wire [63:0] T_158;
  wire [63:0] T_160;
  wire [63:0] T_161;
  wire [61:0] T_165;
  wire [63:0] GEN_25;
  wire [63:0] T_166;
  wire [61:0] T_167;
  wire [63:0] GEN_26;
  wire [63:0] T_168;
  wire [63:0] T_170;
  wire [63:0] T_171;
  wire [62:0] T_175;
  wire [63:0] GEN_27;
  wire [63:0] T_176;
  wire [62:0] T_177;
  wire [63:0] GEN_28;
  wire [63:0] T_178;
  wire [63:0] T_180;
  wire [63:0] shout_l;
  wire [63:0] T_185;
  wire [3:0] GEN_30;
  wire  T_186;
  wire [63:0] T_188;
  wire [63:0] shout;
  wire [3:0] GEN_31;
  wire  T_189;
  wire [3:0] GEN_32;
  wire  T_190;
  wire  T_191;
  wire [63:0] T_193;
  wire [3:0] GEN_34;
  wire  T_195;
  wire  T_196;
  wire [63:0] T_197;
  wire [63:0] T_199;
  wire [63:0] logic$;
  wire [3:0] GEN_35;
  wire  T_200;
  wire [3:0] GEN_36;
  wire  T_201;
  wire  T_202;
  wire  T_203;
  wire  T_204;
  wire  T_205;
  wire [63:0] GEN_37;
  wire [63:0] T_206;
  wire [63:0] shift_logic;
  wire [3:0] GEN_38;
  wire  T_207;
  wire  T_208;
  wire  T_209;
  wire [63:0] out;
  wire  T_213;
  wire  T_214;
  wire [31:0] GEN_39;
  wire [32:0] T_216;
  wire [31:0] T_217;
  wire [31:0] T_218;
  wire [63:0] T_219;
  wire [63:0] GEN_0;
  assign io_out = GEN_0;
  assign io_adder_out = T_13;
  assign io_cmp_out = T_30;
  assign T_7 = io_fn[3];
  assign T_8 = ~ io_in2;
  assign in2_inv = T_7 ? T_8 : io_in2;
  assign in1_xor_in2 = io_in1 ^ in2_inv;
  assign T_9 = io_in1 + in2_inv;
  assign T_10 = T_9[63:0];
  assign GEN_1 = {{63'd0}, T_7};
  assign T_12 = T_10 + GEN_1;
  assign T_13 = T_12[63:0];
  assign T_14 = io_fn[0];
  assign T_17 = T_7 == 1'h0;
  assign GEN_2 = {{63'd0}, 1'h0};
  assign T_19 = in1_xor_in2 == GEN_2;
  assign T_20 = io_in1[63];
  assign T_21 = io_in2[63];
  assign T_22 = T_20 == T_21;
  assign T_23 = io_adder_out[63];
  assign T_24 = io_fn[1];
  assign T_27 = T_24 ? T_21 : T_20;
  assign T_28 = T_22 ? T_23 : T_27;
  assign T_29 = T_17 ? T_19 : T_28;
  assign T_30 = T_14 ^ T_29;
  assign T_32 = io_in1[31];
  assign T_33 = T_7 & T_32;
  assign GEN_3 = {{31'd0}, T_33};
  assign T_35 = 32'h0 - GEN_3;
  assign T_36 = T_35[31:0];
  assign T_41 = io_in1[63:32];
  assign T_42 = io_dw ? T_41 : T_36;
  assign T_43 = io_in2[5];
  assign T_48 = T_43 & io_dw;
  assign T_49 = io_in2[4:0];
  assign shamt = {T_48,T_49};
  assign T_50 = io_in1[31:0];
  assign shin_r = {T_42,T_50};
  assign GEN_4 = {{1'd0}, 3'h5};
  assign T_51 = io_fn == GEN_4;
  assign T_52 = io_fn == 4'hb;
  assign T_53 = T_51 | T_52;
  assign T_58 = shin_r[63:32];
  assign GEN_5 = {{32'd0}, T_58};
  assign T_59 = GEN_5 & 64'hffffffff;
  assign T_60 = shin_r[31:0];
  assign GEN_6 = {{32'd0}, T_60};
  assign T_61 = GEN_6 << 32;
  assign T_63 = T_61 & 64'hffffffff00000000;
  assign T_64 = T_59 | T_63;
  assign T_68 = T_64[63:16];
  assign GEN_7 = {{16'd0}, T_68};
  assign T_69 = GEN_7 & 64'hffff0000ffff;
  assign T_70 = T_64[47:0];
  assign GEN_8 = {{16'd0}, T_70};
  assign T_71 = GEN_8 << 16;
  assign T_73 = T_71 & 64'hffff0000ffff0000;
  assign T_74 = T_69 | T_73;
  assign T_78 = T_74[63:8];
  assign GEN_9 = {{8'd0}, T_78};
  assign T_79 = GEN_9 & 64'hff00ff00ff00ff;
  assign T_80 = T_74[55:0];
  assign GEN_10 = {{8'd0}, T_80};
  assign T_81 = GEN_10 << 8;
  assign T_83 = T_81 & 64'hff00ff00ff00ff00;
  assign T_84 = T_79 | T_83;
  assign T_88 = T_84[63:4];
  assign GEN_11 = {{4'd0}, T_88};
  assign T_89 = GEN_11 & 64'hf0f0f0f0f0f0f0f;
  assign T_90 = T_84[59:0];
  assign GEN_12 = {{4'd0}, T_90};
  assign T_91 = GEN_12 << 4;
  assign T_93 = T_91 & 64'hf0f0f0f0f0f0f0f0;
  assign T_94 = T_89 | T_93;
  assign T_98 = T_94[63:2];
  assign GEN_13 = {{2'd0}, T_98};
  assign T_99 = GEN_13 & 64'h3333333333333333;
  assign T_100 = T_94[61:0];
  assign GEN_14 = {{2'd0}, T_100};
  assign T_101 = GEN_14 << 2;
  assign T_103 = T_101 & 64'hcccccccccccccccc;
  assign T_104 = T_99 | T_103;
  assign T_108 = T_104[63:1];
  assign GEN_15 = {{1'd0}, T_108};
  assign T_109 = GEN_15 & 64'h5555555555555555;
  assign T_110 = T_104[62:0];
  assign GEN_16 = {{1'd0}, T_110};
  assign T_111 = GEN_16 << 1;
  assign T_113 = T_111 & 64'haaaaaaaaaaaaaaaa;
  assign T_114 = T_109 | T_113;
  assign shin = T_53 ? shin_r : T_114;
  assign T_116 = shin[63];
  assign T_117 = T_7 & T_116;
  assign T_118 = {T_117,shin};
  assign T_119 = $signed(T_118);
  assign T_120 = $signed(T_119) >>> shamt;
  assign shout_r = T_120[63:0];
  assign T_125 = shout_r[63:32];
  assign GEN_17 = {{32'd0}, T_125};
  assign T_126 = GEN_17 & 64'hffffffff;
  assign T_127 = shout_r[31:0];
  assign GEN_18 = {{32'd0}, T_127};
  assign T_128 = GEN_18 << 32;
  assign T_130 = T_128 & 64'hffffffff00000000;
  assign T_131 = T_126 | T_130;
  assign T_135 = T_131[63:16];
  assign GEN_19 = {{16'd0}, T_135};
  assign T_136 = GEN_19 & 64'hffff0000ffff;
  assign T_137 = T_131[47:0];
  assign GEN_20 = {{16'd0}, T_137};
  assign T_138 = GEN_20 << 16;
  assign T_140 = T_138 & 64'hffff0000ffff0000;
  assign T_141 = T_136 | T_140;
  assign T_145 = T_141[63:8];
  assign GEN_21 = {{8'd0}, T_145};
  assign T_146 = GEN_21 & 64'hff00ff00ff00ff;
  assign T_147 = T_141[55:0];
  assign GEN_22 = {{8'd0}, T_147};
  assign T_148 = GEN_22 << 8;
  assign T_150 = T_148 & 64'hff00ff00ff00ff00;
  assign T_151 = T_146 | T_150;
  assign T_155 = T_151[63:4];
  assign GEN_23 = {{4'd0}, T_155};
  assign T_156 = GEN_23 & 64'hf0f0f0f0f0f0f0f;
  assign T_157 = T_151[59:0];
  assign GEN_24 = {{4'd0}, T_157};
  assign T_158 = GEN_24 << 4;
  assign T_160 = T_158 & 64'hf0f0f0f0f0f0f0f0;
  assign T_161 = T_156 | T_160;
  assign T_165 = T_161[63:2];
  assign GEN_25 = {{2'd0}, T_165};
  assign T_166 = GEN_25 & 64'h3333333333333333;
  assign T_167 = T_161[61:0];
  assign GEN_26 = {{2'd0}, T_167};
  assign T_168 = GEN_26 << 2;
  assign T_170 = T_168 & 64'hcccccccccccccccc;
  assign T_171 = T_166 | T_170;
  assign T_175 = T_171[63:1];
  assign GEN_27 = {{1'd0}, T_175};
  assign T_176 = GEN_27 & 64'h5555555555555555;
  assign T_177 = T_171[62:0];
  assign GEN_28 = {{1'd0}, T_177};
  assign T_178 = GEN_28 << 1;
  assign T_180 = T_178 & 64'haaaaaaaaaaaaaaaa;
  assign shout_l = T_176 | T_180;
  assign T_185 = T_53 ? shout_r : {{63'd0}, 1'h0};
  assign GEN_30 = {{3'd0}, 1'h1};
  assign T_186 = io_fn == GEN_30;
  assign T_188 = T_186 ? shout_l : {{63'd0}, 1'h0};
  assign shout = T_185 | T_188;
  assign GEN_31 = {{1'd0}, 3'h4};
  assign T_189 = io_fn == GEN_31;
  assign GEN_32 = {{1'd0}, 3'h6};
  assign T_190 = io_fn == GEN_32;
  assign T_191 = T_189 | T_190;
  assign T_193 = T_191 ? in1_xor_in2 : {{63'd0}, 1'h0};
  assign GEN_34 = {{1'd0}, 3'h7};
  assign T_195 = io_fn == GEN_34;
  assign T_196 = T_190 | T_195;
  assign T_197 = io_in1 & io_in2;
  assign T_199 = T_196 ? T_197 : {{63'd0}, 1'h0};
  assign logic$ = T_193 | T_199;
  assign GEN_35 = {{2'd0}, 2'h2};
  assign T_200 = io_fn == GEN_35;
  assign GEN_36 = {{2'd0}, 2'h3};
  assign T_201 = io_fn == GEN_36;
  assign T_202 = T_200 | T_201;
  assign T_203 = io_fn >= 4'hc;
  assign T_204 = T_202 | T_203;
  assign T_205 = T_204 & io_cmp_out;
  assign GEN_37 = {{63'd0}, T_205};
  assign T_206 = GEN_37 | logic$;
  assign shift_logic = T_206 | shout;
  assign GEN_38 = {{3'd0}, 1'h0};
  assign T_207 = io_fn == GEN_38;
  assign T_208 = io_fn == 4'ha;
  assign T_209 = T_207 | T_208;
  assign out = T_209 ? io_adder_out : shift_logic;
  assign T_213 = 1'h0 == io_dw;
  assign T_214 = out[31];
  assign GEN_39 = {{31'd0}, T_214};
  assign T_216 = 32'h0 - GEN_39;
  assign T_217 = T_216[31:0];
  assign T_218 = out[31:0];
  assign T_219 = {T_217,T_218};
  assign GEN_0 = T_213 ? T_219 : out;
endmodule
module MulDiv(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [3:0] io_req_bits_fn,
  input   io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input  [4:0] io_req_bits_tag,
  input   io_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0] io_resp_bits_tag
);
  reg [2:0] state;
  reg [31:0] GEN_43;
  reg [3:0] req_fn;
  reg [31:0] GEN_44;
  reg  req_dw;
  reg [31:0] GEN_47;
  reg [63:0] req_in1;
  reg [63:0] GEN_48;
  reg [63:0] req_in2;
  reg [63:0] GEN_49;
  reg [4:0] req_tag;
  reg [31:0] GEN_52;
  reg [6:0] count;
  reg [31:0] GEN_54;
  reg  neg_out;
  reg [31:0] GEN_55;
  reg  isMul;
  reg [31:0] GEN_56;
  reg  isHi;
  reg [31:0] GEN_57;
  reg [64:0] divisor;
  reg [95:0] GEN_58;
  reg [129:0] remainder;
  reg [159:0] GEN_59;
  wire [3:0] T_62;
  wire  T_64;
  wire [3:0] T_66;
  wire  T_68;
  wire  T_71;
  wire [3:0] T_73;
  wire  T_75;
  wire [3:0] T_77;
  wire  T_79;
  wire  T_82;
  wire  T_83;
  wire [3:0] T_85;
  wire  T_87;
  wire [3:0] T_89;
  wire  T_91;
  wire  T_94;
  wire  T_95;
  wire  T_103;
  wire  T_105;
  wire  T_106;
  wire  T_107;
  wire  lhs_sign;
  wire [31:0] GEN_34;
  wire [32:0] T_109;
  wire [31:0] T_110;
  wire [31:0] T_111;
  wire [31:0] T_112;
  wire [31:0] T_113;
  wire [63:0] lhs_in;
  wire  T_120;
  wire  T_121;
  wire  T_122;
  wire  rhs_sign;
  wire [31:0] GEN_35;
  wire [32:0] T_124;
  wire [31:0] T_125;
  wire [31:0] T_126;
  wire [31:0] T_127;
  wire [31:0] T_128;
  wire [63:0] rhs_in;
  wire [64:0] T_129;
  wire [65:0] T_131;
  wire [64:0] subtractor;
  wire  less;
  wire [63:0] T_132;
  wire [63:0] GEN_36;
  wire [64:0] T_134;
  wire [63:0] negated_remainder;
  wire  T_135;
  wire  T_136;
  wire  T_137;
  wire [129:0] GEN_0;
  wire  T_138;
  wire  T_139;
  wire [64:0] GEN_1;
  wire [129:0] GEN_2;
  wire [64:0] GEN_3;
  wire [2:0] GEN_4;
  wire  T_140;
  wire [129:0] GEN_5;
  wire [2:0] GEN_6;
  wire  T_141;
  wire [63:0] T_142;
  wire [2:0] T_143;
  wire [129:0] GEN_7;
  wire [2:0] GEN_8;
  wire  T_144;
  wire  T_145;
  wire [64:0] T_146;
  wire [128:0] T_148;
  wire [63:0] T_149;
  wire [64:0] T_150;
  wire [64:0] T_151;
  wire [64:0] T_152;
  wire [7:0] T_153;
  wire [64:0] GEN_37;
  wire [72:0] T_154;
  wire [72:0] GEN_38;
  wire [73:0] T_155;
  wire [72:0] T_156;
  wire [72:0] T_157;
  wire [55:0] T_158;
  wire [72:0] T_159;
  wire [128:0] T_160;
  wire [6:0] GEN_39;
  wire [10:0] T_163;
  wire [5:0] T_164;
  wire [64:0] GEN_40;
  wire [64:0] T_165;
  wire [63:0] T_166;
  wire [6:0] GEN_41;
  wire  T_169;
  wire [6:0] GEN_42;
  wire  T_172;
  wire  T_173;
  wire  T_175;
  wire  T_176;
  wire [63:0] T_177;
  wire [63:0] T_178;
  wire  T_180;
  wire  T_181;
  wire [10:0] GEN_45;
  wire [11:0] T_185;
  wire [10:0] T_186;
  wire [5:0] T_187;
  wire [128:0] T_188;
  wire [64:0] T_189;
  wire [128:0] T_190;
  wire [63:0] T_191;
  wire [128:0] T_192;
  wire [64:0] T_193;
  wire [63:0] T_195;
  wire [65:0] T_196;
  wire [129:0] T_197;
  wire [6:0] GEN_46;
  wire [7:0] T_199;
  wire [6:0] T_200;
  wire  T_202;
  wire  T_203;
  wire [2:0] T_204;
  wire [2:0] GEN_9;
  wire [129:0] GEN_10;
  wire [6:0] GEN_11;
  wire [2:0] GEN_12;
  wire  T_207;
  wire  T_208;
  wire  T_210;
  wire [2:0] T_212;
  wire [2:0] GEN_13;
  wire [63:0] T_216;
  wire [63:0] T_217;
  wire [63:0] T_218;
  wire  T_221;
  wire [127:0] T_222;
  wire [128:0] T_223;
  wire [63:0] T_224;
  wire  T_225;
  wire  T_227;
  wire  T_229;
  wire  T_231;
  wire  T_233;
  wire  T_235;
  wire  T_237;
  wire  T_239;
  wire  T_241;
  wire  T_243;
  wire  T_245;
  wire  T_247;
  wire  T_249;
  wire  T_251;
  wire  T_253;
  wire  T_255;
  wire  T_257;
  wire  T_259;
  wire  T_261;
  wire  T_263;
  wire  T_265;
  wire  T_267;
  wire  T_269;
  wire  T_271;
  wire  T_273;
  wire  T_275;
  wire  T_277;
  wire  T_279;
  wire  T_281;
  wire  T_283;
  wire  T_285;
  wire  T_287;
  wire  T_289;
  wire  T_291;
  wire  T_293;
  wire  T_295;
  wire  T_297;
  wire  T_299;
  wire  T_301;
  wire  T_303;
  wire  T_305;
  wire  T_307;
  wire  T_309;
  wire  T_311;
  wire  T_313;
  wire  T_315;
  wire  T_317;
  wire  T_319;
  wire  T_321;
  wire  T_323;
  wire  T_325;
  wire  T_327;
  wire  T_329;
  wire  T_331;
  wire  T_333;
  wire  T_335;
  wire  T_337;
  wire  T_339;
  wire  T_341;
  wire  T_343;
  wire  T_345;
  wire  T_347;
  wire  T_349;
  wire [1:0] T_351;
  wire [1:0] T_352;
  wire [2:0] T_353;
  wire [2:0] T_354;
  wire [2:0] T_355;
  wire [2:0] T_356;
  wire [3:0] T_357;
  wire [3:0] T_358;
  wire [3:0] T_359;
  wire [3:0] T_360;
  wire [3:0] T_361;
  wire [3:0] T_362;
  wire [3:0] T_363;
  wire [3:0] T_364;
  wire [4:0] T_365;
  wire [4:0] T_366;
  wire [4:0] T_367;
  wire [4:0] T_368;
  wire [4:0] T_369;
  wire [4:0] T_370;
  wire [4:0] T_371;
  wire [4:0] T_372;
  wire [4:0] T_373;
  wire [4:0] T_374;
  wire [4:0] T_375;
  wire [4:0] T_376;
  wire [4:0] T_377;
  wire [4:0] T_378;
  wire [4:0] T_379;
  wire [4:0] T_380;
  wire [5:0] T_381;
  wire [5:0] T_382;
  wire [5:0] T_383;
  wire [5:0] T_384;
  wire [5:0] T_385;
  wire [5:0] T_386;
  wire [5:0] T_387;
  wire [5:0] T_388;
  wire [5:0] T_389;
  wire [5:0] T_390;
  wire [5:0] T_391;
  wire [5:0] T_392;
  wire [5:0] T_393;
  wire [5:0] T_394;
  wire [5:0] T_395;
  wire [5:0] T_396;
  wire [5:0] T_397;
  wire [5:0] T_398;
  wire [5:0] T_399;
  wire [5:0] T_400;
  wire [5:0] T_401;
  wire [5:0] T_402;
  wire [5:0] T_403;
  wire [5:0] T_404;
  wire [5:0] T_405;
  wire [5:0] T_406;
  wire [5:0] T_407;
  wire [5:0] T_408;
  wire [5:0] T_409;
  wire [5:0] T_410;
  wire [5:0] T_411;
  wire [5:0] T_412;
  wire  T_414;
  wire  T_416;
  wire  T_418;
  wire  T_420;
  wire  T_422;
  wire  T_424;
  wire  T_426;
  wire  T_428;
  wire  T_430;
  wire  T_432;
  wire  T_434;
  wire  T_436;
  wire  T_438;
  wire  T_440;
  wire  T_442;
  wire  T_444;
  wire  T_446;
  wire  T_448;
  wire  T_450;
  wire  T_452;
  wire  T_454;
  wire  T_456;
  wire  T_458;
  wire  T_460;
  wire  T_462;
  wire  T_464;
  wire  T_466;
  wire  T_468;
  wire  T_470;
  wire  T_472;
  wire  T_474;
  wire  T_476;
  wire  T_478;
  wire  T_480;
  wire  T_482;
  wire  T_484;
  wire  T_486;
  wire  T_488;
  wire  T_490;
  wire  T_492;
  wire  T_494;
  wire  T_496;
  wire  T_498;
  wire  T_500;
  wire  T_502;
  wire  T_504;
  wire  T_506;
  wire  T_508;
  wire  T_510;
  wire  T_512;
  wire  T_514;
  wire  T_516;
  wire  T_518;
  wire  T_520;
  wire  T_522;
  wire  T_524;
  wire  T_526;
  wire  T_528;
  wire  T_530;
  wire  T_532;
  wire  T_534;
  wire  T_536;
  wire  T_538;
  wire [1:0] T_540;
  wire [1:0] T_541;
  wire [2:0] T_542;
  wire [2:0] T_543;
  wire [2:0] T_544;
  wire [2:0] T_545;
  wire [3:0] T_546;
  wire [3:0] T_547;
  wire [3:0] T_548;
  wire [3:0] T_549;
  wire [3:0] T_550;
  wire [3:0] T_551;
  wire [3:0] T_552;
  wire [3:0] T_553;
  wire [4:0] T_554;
  wire [4:0] T_555;
  wire [4:0] T_556;
  wire [4:0] T_557;
  wire [4:0] T_558;
  wire [4:0] T_559;
  wire [4:0] T_560;
  wire [4:0] T_561;
  wire [4:0] T_562;
  wire [4:0] T_563;
  wire [4:0] T_564;
  wire [4:0] T_565;
  wire [4:0] T_566;
  wire [4:0] T_567;
  wire [4:0] T_568;
  wire [4:0] T_569;
  wire [5:0] T_570;
  wire [5:0] T_571;
  wire [5:0] T_572;
  wire [5:0] T_573;
  wire [5:0] T_574;
  wire [5:0] T_575;
  wire [5:0] T_576;
  wire [5:0] T_577;
  wire [5:0] T_578;
  wire [5:0] T_579;
  wire [5:0] T_580;
  wire [5:0] T_581;
  wire [5:0] T_582;
  wire [5:0] T_583;
  wire [5:0] T_584;
  wire [5:0] T_585;
  wire [5:0] T_586;
  wire [5:0] T_587;
  wire [5:0] T_588;
  wire [5:0] T_589;
  wire [5:0] T_590;
  wire [5:0] T_591;
  wire [5:0] T_592;
  wire [5:0] T_593;
  wire [5:0] T_594;
  wire [5:0] T_595;
  wire [5:0] T_596;
  wire [5:0] T_597;
  wire [5:0] T_598;
  wire [5:0] T_599;
  wire [5:0] T_600;
  wire [5:0] T_601;
  wire [6:0] T_603;
  wire [5:0] T_604;
  wire [6:0] T_605;
  wire [5:0] T_606;
  wire  T_607;
  wire  T_609;
  wire  T_610;
  wire [5:0] GEN_50;
  wire  T_612;
  wire  T_613;
  wire  T_614;
  wire [5:0] T_619;
  wire [126:0] GEN_51;
  wire [126:0] T_621;
  wire [128:0] GEN_14;
  wire [6:0] GEN_15;
  wire  T_626;
  wire  T_629;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [6:0] GEN_18;
  wire [129:0] GEN_19;
  wire  GEN_20;
  wire  T_631;
  wire  T_632;
  wire [2:0] GEN_21;
  wire  T_633;
  wire  T_635;
  wire  T_636;
  wire  T_637;
  wire [2:0] T_638;
  wire  T_642;
  wire  T_643;
  wire  T_644;
  wire [64:0] T_645;
  wire [2:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [6:0] GEN_25;
  wire  GEN_26;
  wire [64:0] GEN_27;
  wire [129:0] GEN_28;
  wire [3:0] GEN_29;
  wire  GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [4:0] GEN_33;
  wire  T_650;
  wire  T_652;
  wire [31:0] GEN_53;
  wire [32:0] T_654;
  wire [31:0] T_655;
  wire [31:0] T_656;
  wire [63:0] T_657;
  wire [63:0] T_659;
  wire  T_660;
  wire  T_661;
  assign io_req_ready = T_661;
  assign io_resp_valid = T_660;
  assign io_resp_bits_data = T_659;
  assign io_resp_bits_tag = req_tag;
  assign T_62 = io_req_bits_fn & 4'h4;
  assign T_64 = T_62 == 4'h0;
  assign T_66 = io_req_bits_fn & 4'h8;
  assign T_68 = T_66 == 4'h8;
  assign T_71 = T_64 | T_68;
  assign T_73 = io_req_bits_fn & 4'h5;
  assign T_75 = T_73 == 4'h1;
  assign T_77 = io_req_bits_fn & 4'h2;
  assign T_79 = T_77 == 4'h2;
  assign T_82 = T_75 | T_79;
  assign T_83 = T_82 | T_68;
  assign T_85 = io_req_bits_fn & 4'h9;
  assign T_87 = T_85 == 4'h0;
  assign T_89 = io_req_bits_fn & 4'h3;
  assign T_91 = T_89 == 4'h0;
  assign T_94 = T_87 | T_64;
  assign T_95 = T_94 | T_91;
  assign T_103 = 1'h0 == io_req_bits_dw;
  assign T_105 = io_req_bits_in1[31];
  assign T_106 = io_req_bits_in1[63];
  assign T_107 = T_103 ? T_105 : T_106;
  assign lhs_sign = T_95 & T_107;
  assign GEN_34 = {{31'd0}, lhs_sign};
  assign T_109 = 32'h0 - GEN_34;
  assign T_110 = T_109[31:0];
  assign T_111 = io_req_bits_in1[63:32];
  assign T_112 = T_103 ? T_110 : T_111;
  assign T_113 = io_req_bits_in1[31:0];
  assign lhs_in = {T_112,T_113};
  assign T_120 = io_req_bits_in2[31];
  assign T_121 = io_req_bits_in2[63];
  assign T_122 = T_103 ? T_120 : T_121;
  assign rhs_sign = T_94 & T_122;
  assign GEN_35 = {{31'd0}, rhs_sign};
  assign T_124 = 32'h0 - GEN_35;
  assign T_125 = T_124[31:0];
  assign T_126 = io_req_bits_in2[63:32];
  assign T_127 = T_103 ? T_125 : T_126;
  assign T_128 = io_req_bits_in2[31:0];
  assign rhs_in = {T_127,T_128};
  assign T_129 = remainder[128:64];
  assign T_131 = T_129 - divisor;
  assign subtractor = T_131[64:0];
  assign less = subtractor[64];
  assign T_132 = remainder[63:0];
  assign GEN_36 = {{63'd0}, 1'h0};
  assign T_134 = GEN_36 - T_132;
  assign negated_remainder = T_134[63:0];
  assign T_135 = state == 3'h1;
  assign T_136 = remainder[63];
  assign T_137 = T_136 | isMul;
  assign GEN_0 = T_137 ? {{66'd0}, negated_remainder} : remainder;
  assign T_138 = divisor[63];
  assign T_139 = T_138 | isMul;
  assign GEN_1 = T_139 ? subtractor : divisor;
  assign GEN_2 = T_135 ? GEN_0 : remainder;
  assign GEN_3 = T_135 ? GEN_1 : divisor;
  assign GEN_4 = T_135 ? 3'h2 : state;
  assign T_140 = state == 3'h4;
  assign GEN_5 = T_140 ? {{66'd0}, negated_remainder} : GEN_2;
  assign GEN_6 = T_140 ? 3'h5 : GEN_4;
  assign T_141 = state == 3'h3;
  assign T_142 = remainder[128:65];
  assign T_143 = neg_out ? 3'h4 : 3'h5;
  assign GEN_7 = T_141 ? {{66'd0}, T_142} : GEN_5;
  assign GEN_8 = T_141 ? T_143 : GEN_6;
  assign T_144 = state == 3'h2;
  assign T_145 = T_144 & isMul;
  assign T_146 = remainder[129:65];
  assign T_148 = {T_146,T_132};
  assign T_149 = T_148[63:0];
  assign T_150 = T_148[128:64];
  assign T_151 = $signed(T_150);
  assign T_152 = $signed(divisor);
  assign T_153 = T_149[7:0];
  assign GEN_37 = {{57'd0}, T_153};
  assign T_154 = $signed(T_152) * $signed({1'b0,GEN_37});
  assign GEN_38 = {{8{T_151[64]}},T_151};
  assign T_155 = $signed(T_154) + $signed(GEN_38);
  assign T_156 = T_155[72:0];
  assign T_157 = $signed(T_156);
  assign T_158 = T_149[63:8];
  assign T_159 = $unsigned(T_157);
  assign T_160 = {T_159,T_158};
  assign GEN_39 = {{3'd0}, 4'h8};
  assign T_163 = count * GEN_39;
  assign T_164 = T_163[5:0];
  assign GEN_40 = $signed(65'h10000000000000000);
  assign T_165 = $signed(GEN_40) >>> T_164;
  assign T_166 = T_165[63:0];
  assign GEN_41 = {{4'd0}, 3'h7};
  assign T_169 = count != GEN_41;
  assign GEN_42 = {{6'd0}, 1'h0};
  assign T_172 = count != GEN_42;
  assign T_173 = T_169 & T_172;
  assign T_175 = isHi == 1'h0;
  assign T_176 = T_173 & T_175;
  assign T_177 = ~ T_166;
  assign T_178 = T_149 & T_177;
  assign T_180 = T_178 == GEN_36;
  assign T_181 = T_176 & T_180;
  assign GEN_45 = {{4'd0}, 7'h40};
  assign T_185 = GEN_45 - T_163;
  assign T_186 = T_185[10:0];
  assign T_187 = T_186[5:0];
  assign T_188 = T_148 >> T_187;
  assign T_189 = T_160[128:64];
  assign T_190 = T_181 ? T_188 : T_160;
  assign T_191 = T_190[63:0];
  assign T_192 = {T_189,T_191};
  assign T_193 = T_192[128:64];
  assign T_195 = T_192[63:0];
  assign T_196 = {T_193,1'h0};
  assign T_197 = {T_196,T_195};
  assign GEN_46 = {{6'd0}, 1'h1};
  assign T_199 = count + GEN_46;
  assign T_200 = T_199[6:0];
  assign T_202 = count == GEN_41;
  assign T_203 = T_181 | T_202;
  assign T_204 = isHi ? 3'h3 : 3'h5;
  assign GEN_9 = T_203 ? T_204 : GEN_8;
  assign GEN_10 = T_145 ? T_197 : GEN_7;
  assign GEN_11 = T_145 ? T_200 : count;
  assign GEN_12 = T_145 ? GEN_9 : GEN_8;
  assign T_207 = isMul == 1'h0;
  assign T_208 = T_144 & T_207;
  assign T_210 = count == 7'h40;
  assign T_212 = isHi ? 3'h3 : T_143;
  assign GEN_13 = T_210 ? T_212 : GEN_12;
  assign T_216 = remainder[127:64];
  assign T_217 = subtractor[63:0];
  assign T_218 = less ? T_216 : T_217;
  assign T_221 = less == 1'h0;
  assign T_222 = {T_218,T_132};
  assign T_223 = {T_222,T_221};
  assign T_224 = divisor[63:0];
  assign T_225 = T_224[63];
  assign T_227 = T_224[62];
  assign T_229 = T_224[61];
  assign T_231 = T_224[60];
  assign T_233 = T_224[59];
  assign T_235 = T_224[58];
  assign T_237 = T_224[57];
  assign T_239 = T_224[56];
  assign T_241 = T_224[55];
  assign T_243 = T_224[54];
  assign T_245 = T_224[53];
  assign T_247 = T_224[52];
  assign T_249 = T_224[51];
  assign T_251 = T_224[50];
  assign T_253 = T_224[49];
  assign T_255 = T_224[48];
  assign T_257 = T_224[47];
  assign T_259 = T_224[46];
  assign T_261 = T_224[45];
  assign T_263 = T_224[44];
  assign T_265 = T_224[43];
  assign T_267 = T_224[42];
  assign T_269 = T_224[41];
  assign T_271 = T_224[40];
  assign T_273 = T_224[39];
  assign T_275 = T_224[38];
  assign T_277 = T_224[37];
  assign T_279 = T_224[36];
  assign T_281 = T_224[35];
  assign T_283 = T_224[34];
  assign T_285 = T_224[33];
  assign T_287 = T_224[32];
  assign T_289 = T_224[31];
  assign T_291 = T_224[30];
  assign T_293 = T_224[29];
  assign T_295 = T_224[28];
  assign T_297 = T_224[27];
  assign T_299 = T_224[26];
  assign T_301 = T_224[25];
  assign T_303 = T_224[24];
  assign T_305 = T_224[23];
  assign T_307 = T_224[22];
  assign T_309 = T_224[21];
  assign T_311 = T_224[20];
  assign T_313 = T_224[19];
  assign T_315 = T_224[18];
  assign T_317 = T_224[17];
  assign T_319 = T_224[16];
  assign T_321 = T_224[15];
  assign T_323 = T_224[14];
  assign T_325 = T_224[13];
  assign T_327 = T_224[12];
  assign T_329 = T_224[11];
  assign T_331 = T_224[10];
  assign T_333 = T_224[9];
  assign T_335 = T_224[8];
  assign T_337 = T_224[7];
  assign T_339 = T_224[6];
  assign T_341 = T_224[5];
  assign T_343 = T_224[4];
  assign T_345 = T_224[3];
  assign T_347 = T_224[2];
  assign T_349 = T_224[1];
  assign T_351 = T_347 ? 2'h2 : {{1'd0}, T_349};
  assign T_352 = T_345 ? 2'h3 : T_351;
  assign T_353 = T_343 ? 3'h4 : {{1'd0}, T_352};
  assign T_354 = T_341 ? 3'h5 : T_353;
  assign T_355 = T_339 ? 3'h6 : T_354;
  assign T_356 = T_337 ? 3'h7 : T_355;
  assign T_357 = T_335 ? 4'h8 : {{1'd0}, T_356};
  assign T_358 = T_333 ? 4'h9 : T_357;
  assign T_359 = T_331 ? 4'ha : T_358;
  assign T_360 = T_329 ? 4'hb : T_359;
  assign T_361 = T_327 ? 4'hc : T_360;
  assign T_362 = T_325 ? 4'hd : T_361;
  assign T_363 = T_323 ? 4'he : T_362;
  assign T_364 = T_321 ? 4'hf : T_363;
  assign T_365 = T_319 ? 5'h10 : {{1'd0}, T_364};
  assign T_366 = T_317 ? 5'h11 : T_365;
  assign T_367 = T_315 ? 5'h12 : T_366;
  assign T_368 = T_313 ? 5'h13 : T_367;
  assign T_369 = T_311 ? 5'h14 : T_368;
  assign T_370 = T_309 ? 5'h15 : T_369;
  assign T_371 = T_307 ? 5'h16 : T_370;
  assign T_372 = T_305 ? 5'h17 : T_371;
  assign T_373 = T_303 ? 5'h18 : T_372;
  assign T_374 = T_301 ? 5'h19 : T_373;
  assign T_375 = T_299 ? 5'h1a : T_374;
  assign T_376 = T_297 ? 5'h1b : T_375;
  assign T_377 = T_295 ? 5'h1c : T_376;
  assign T_378 = T_293 ? 5'h1d : T_377;
  assign T_379 = T_291 ? 5'h1e : T_378;
  assign T_380 = T_289 ? 5'h1f : T_379;
  assign T_381 = T_287 ? 6'h20 : {{1'd0}, T_380};
  assign T_382 = T_285 ? 6'h21 : T_381;
  assign T_383 = T_283 ? 6'h22 : T_382;
  assign T_384 = T_281 ? 6'h23 : T_383;
  assign T_385 = T_279 ? 6'h24 : T_384;
  assign T_386 = T_277 ? 6'h25 : T_385;
  assign T_387 = T_275 ? 6'h26 : T_386;
  assign T_388 = T_273 ? 6'h27 : T_387;
  assign T_389 = T_271 ? 6'h28 : T_388;
  assign T_390 = T_269 ? 6'h29 : T_389;
  assign T_391 = T_267 ? 6'h2a : T_390;
  assign T_392 = T_265 ? 6'h2b : T_391;
  assign T_393 = T_263 ? 6'h2c : T_392;
  assign T_394 = T_261 ? 6'h2d : T_393;
  assign T_395 = T_259 ? 6'h2e : T_394;
  assign T_396 = T_257 ? 6'h2f : T_395;
  assign T_397 = T_255 ? 6'h30 : T_396;
  assign T_398 = T_253 ? 6'h31 : T_397;
  assign T_399 = T_251 ? 6'h32 : T_398;
  assign T_400 = T_249 ? 6'h33 : T_399;
  assign T_401 = T_247 ? 6'h34 : T_400;
  assign T_402 = T_245 ? 6'h35 : T_401;
  assign T_403 = T_243 ? 6'h36 : T_402;
  assign T_404 = T_241 ? 6'h37 : T_403;
  assign T_405 = T_239 ? 6'h38 : T_404;
  assign T_406 = T_237 ? 6'h39 : T_405;
  assign T_407 = T_235 ? 6'h3a : T_406;
  assign T_408 = T_233 ? 6'h3b : T_407;
  assign T_409 = T_231 ? 6'h3c : T_408;
  assign T_410 = T_229 ? 6'h3d : T_409;
  assign T_411 = T_227 ? 6'h3e : T_410;
  assign T_412 = T_225 ? 6'h3f : T_411;
  assign T_414 = T_132[63];
  assign T_416 = T_132[62];
  assign T_418 = T_132[61];
  assign T_420 = T_132[60];
  assign T_422 = T_132[59];
  assign T_424 = T_132[58];
  assign T_426 = T_132[57];
  assign T_428 = T_132[56];
  assign T_430 = T_132[55];
  assign T_432 = T_132[54];
  assign T_434 = T_132[53];
  assign T_436 = T_132[52];
  assign T_438 = T_132[51];
  assign T_440 = T_132[50];
  assign T_442 = T_132[49];
  assign T_444 = T_132[48];
  assign T_446 = T_132[47];
  assign T_448 = T_132[46];
  assign T_450 = T_132[45];
  assign T_452 = T_132[44];
  assign T_454 = T_132[43];
  assign T_456 = T_132[42];
  assign T_458 = T_132[41];
  assign T_460 = T_132[40];
  assign T_462 = T_132[39];
  assign T_464 = T_132[38];
  assign T_466 = T_132[37];
  assign T_468 = T_132[36];
  assign T_470 = T_132[35];
  assign T_472 = T_132[34];
  assign T_474 = T_132[33];
  assign T_476 = T_132[32];
  assign T_478 = T_132[31];
  assign T_480 = T_132[30];
  assign T_482 = T_132[29];
  assign T_484 = T_132[28];
  assign T_486 = T_132[27];
  assign T_488 = T_132[26];
  assign T_490 = T_132[25];
  assign T_492 = T_132[24];
  assign T_494 = T_132[23];
  assign T_496 = T_132[22];
  assign T_498 = T_132[21];
  assign T_500 = T_132[20];
  assign T_502 = T_132[19];
  assign T_504 = T_132[18];
  assign T_506 = T_132[17];
  assign T_508 = T_132[16];
  assign T_510 = T_132[15];
  assign T_512 = T_132[14];
  assign T_514 = T_132[13];
  assign T_516 = T_132[12];
  assign T_518 = T_132[11];
  assign T_520 = T_132[10];
  assign T_522 = T_132[9];
  assign T_524 = T_132[8];
  assign T_526 = T_132[7];
  assign T_528 = T_132[6];
  assign T_530 = T_132[5];
  assign T_532 = T_132[4];
  assign T_534 = T_132[3];
  assign T_536 = T_132[2];
  assign T_538 = T_132[1];
  assign T_540 = T_536 ? 2'h2 : {{1'd0}, T_538};
  assign T_541 = T_534 ? 2'h3 : T_540;
  assign T_542 = T_532 ? 3'h4 : {{1'd0}, T_541};
  assign T_543 = T_530 ? 3'h5 : T_542;
  assign T_544 = T_528 ? 3'h6 : T_543;
  assign T_545 = T_526 ? 3'h7 : T_544;
  assign T_546 = T_524 ? 4'h8 : {{1'd0}, T_545};
  assign T_547 = T_522 ? 4'h9 : T_546;
  assign T_548 = T_520 ? 4'ha : T_547;
  assign T_549 = T_518 ? 4'hb : T_548;
  assign T_550 = T_516 ? 4'hc : T_549;
  assign T_551 = T_514 ? 4'hd : T_550;
  assign T_552 = T_512 ? 4'he : T_551;
  assign T_553 = T_510 ? 4'hf : T_552;
  assign T_554 = T_508 ? 5'h10 : {{1'd0}, T_553};
  assign T_555 = T_506 ? 5'h11 : T_554;
  assign T_556 = T_504 ? 5'h12 : T_555;
  assign T_557 = T_502 ? 5'h13 : T_556;
  assign T_558 = T_500 ? 5'h14 : T_557;
  assign T_559 = T_498 ? 5'h15 : T_558;
  assign T_560 = T_496 ? 5'h16 : T_559;
  assign T_561 = T_494 ? 5'h17 : T_560;
  assign T_562 = T_492 ? 5'h18 : T_561;
  assign T_563 = T_490 ? 5'h19 : T_562;
  assign T_564 = T_488 ? 5'h1a : T_563;
  assign T_565 = T_486 ? 5'h1b : T_564;
  assign T_566 = T_484 ? 5'h1c : T_565;
  assign T_567 = T_482 ? 5'h1d : T_566;
  assign T_568 = T_480 ? 5'h1e : T_567;
  assign T_569 = T_478 ? 5'h1f : T_568;
  assign T_570 = T_476 ? 6'h20 : {{1'd0}, T_569};
  assign T_571 = T_474 ? 6'h21 : T_570;
  assign T_572 = T_472 ? 6'h22 : T_571;
  assign T_573 = T_470 ? 6'h23 : T_572;
  assign T_574 = T_468 ? 6'h24 : T_573;
  assign T_575 = T_466 ? 6'h25 : T_574;
  assign T_576 = T_464 ? 6'h26 : T_575;
  assign T_577 = T_462 ? 6'h27 : T_576;
  assign T_578 = T_460 ? 6'h28 : T_577;
  assign T_579 = T_458 ? 6'h29 : T_578;
  assign T_580 = T_456 ? 6'h2a : T_579;
  assign T_581 = T_454 ? 6'h2b : T_580;
  assign T_582 = T_452 ? 6'h2c : T_581;
  assign T_583 = T_450 ? 6'h2d : T_582;
  assign T_584 = T_448 ? 6'h2e : T_583;
  assign T_585 = T_446 ? 6'h2f : T_584;
  assign T_586 = T_444 ? 6'h30 : T_585;
  assign T_587 = T_442 ? 6'h31 : T_586;
  assign T_588 = T_440 ? 6'h32 : T_587;
  assign T_589 = T_438 ? 6'h33 : T_588;
  assign T_590 = T_436 ? 6'h34 : T_589;
  assign T_591 = T_434 ? 6'h35 : T_590;
  assign T_592 = T_432 ? 6'h36 : T_591;
  assign T_593 = T_430 ? 6'h37 : T_592;
  assign T_594 = T_428 ? 6'h38 : T_593;
  assign T_595 = T_426 ? 6'h39 : T_594;
  assign T_596 = T_424 ? 6'h3a : T_595;
  assign T_597 = T_422 ? 6'h3b : T_596;
  assign T_598 = T_420 ? 6'h3c : T_597;
  assign T_599 = T_418 ? 6'h3d : T_598;
  assign T_600 = T_416 ? 6'h3e : T_599;
  assign T_601 = T_414 ? 6'h3f : T_600;
  assign T_603 = 6'h3f + T_412;
  assign T_604 = T_603[5:0];
  assign T_605 = T_604 - T_601;
  assign T_606 = T_605[5:0];
  assign T_607 = T_412 > T_601;
  assign T_609 = count == GEN_42;
  assign T_610 = T_609 & less;
  assign GEN_50 = {{5'd0}, 1'h0};
  assign T_612 = T_606 > GEN_50;
  assign T_613 = T_612 | T_607;
  assign T_614 = T_610 & T_613;
  assign T_619 = T_607 ? 6'h3f : T_606;
  assign GEN_51 = {{63'd0}, T_132};
  assign T_621 = GEN_51 << T_619;
  assign GEN_14 = T_614 ? {{2'd0}, T_621} : T_223;
  assign GEN_15 = T_614 ? {{1'd0}, T_619} : T_200;
  assign T_626 = T_609 & T_221;
  assign T_629 = T_626 & T_175;
  assign GEN_16 = T_629 ? 1'h0 : neg_out;
  assign GEN_17 = T_208 ? GEN_13 : GEN_12;
  assign GEN_18 = T_208 ? GEN_15 : GEN_11;
  assign GEN_19 = T_208 ? {{1'd0}, GEN_14} : GEN_10;
  assign GEN_20 = T_208 ? GEN_16 : neg_out;
  assign T_631 = io_resp_ready & io_resp_valid;
  assign T_632 = T_631 | io_kill;
  assign GEN_21 = T_632 ? 3'h0 : GEN_17;
  assign T_633 = io_req_ready & io_req_valid;
  assign T_635 = T_71 == 1'h0;
  assign T_636 = rhs_sign & T_635;
  assign T_637 = lhs_sign | T_636;
  assign T_638 = T_637 ? 3'h1 : 3'h2;
  assign T_642 = lhs_sign != rhs_sign;
  assign T_643 = T_83 ? lhs_sign : T_642;
  assign T_644 = T_635 & T_643;
  assign T_645 = {rhs_sign,rhs_in};
  assign GEN_22 = T_633 ? T_638 : GEN_21;
  assign GEN_23 = T_633 ? T_71 : isMul;
  assign GEN_24 = T_633 ? T_83 : isHi;
  assign GEN_25 = T_633 ? {{6'd0}, 1'h0} : GEN_18;
  assign GEN_26 = T_633 ? T_644 : GEN_20;
  assign GEN_27 = T_633 ? T_645 : GEN_3;
  assign GEN_28 = T_633 ? {{66'd0}, lhs_in} : GEN_19;
  assign GEN_29 = T_633 ? io_req_bits_fn : req_fn;
  assign GEN_30 = T_633 ? io_req_bits_dw : req_dw;
  assign GEN_31 = T_633 ? io_req_bits_in1 : req_in1;
  assign GEN_32 = T_633 ? io_req_bits_in2 : req_in2;
  assign GEN_33 = T_633 ? io_req_bits_tag : req_tag;
  assign T_650 = 1'h0 == req_dw;
  assign T_652 = remainder[31];
  assign GEN_53 = {{31'd0}, T_652};
  assign T_654 = 32'h0 - GEN_53;
  assign T_655 = T_654[31:0];
  assign T_656 = remainder[31:0];
  assign T_657 = {T_655,T_656};
  assign T_659 = T_650 ? T_657 : T_132;
  assign T_660 = state == 3'h5;
  assign T_661 = state == 3'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_43 = {1{$random}};
  state = GEN_43[2:0];
  GEN_44 = {1{$random}};
  req_fn = GEN_44[3:0];
  GEN_47 = {1{$random}};
  req_dw = GEN_47[0:0];
  GEN_48 = {2{$random}};
  req_in1 = GEN_48[63:0];
  GEN_49 = {2{$random}};
  req_in2 = GEN_49[63:0];
  GEN_52 = {1{$random}};
  req_tag = GEN_52[4:0];
  GEN_54 = {1{$random}};
  count = GEN_54[6:0];
  GEN_55 = {1{$random}};
  neg_out = GEN_55[0:0];
  GEN_56 = {1{$random}};
  isMul = GEN_56[0:0];
  GEN_57 = {1{$random}};
  isHi = GEN_57[0:0];
  GEN_58 = {3{$random}};
  divisor = GEN_58[64:0];
  GEN_59 = {5{$random}};
  remainder = GEN_59[129:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      if(T_633) begin
        if(T_637) begin
          state <= 3'h1;
        end else begin
          state <= 3'h2;
        end
      end else begin
        if(T_632) begin
          state <= 3'h0;
        end else begin
          if(T_208) begin
            if(T_210) begin
              if(isHi) begin
                state <= 3'h3;
              end else begin
                if(neg_out) begin
                  state <= 3'h4;
                end else begin
                  state <= 3'h5;
                end
              end
            end else begin
              if(T_145) begin
                if(T_203) begin
                  if(isHi) begin
                    state <= 3'h3;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_141) begin
                    if(neg_out) begin
                      state <= 3'h4;
                    end else begin
                      state <= 3'h5;
                    end
                  end else begin
                    if(T_140) begin
                      state <= 3'h5;
                    end else begin
                      if(T_135) begin
                        state <= 3'h2;
                      end
                    end
                  end
                end
              end else begin
                if(T_141) begin
                  if(neg_out) begin
                    state <= 3'h4;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_140) begin
                    state <= 3'h5;
                  end else begin
                    if(T_135) begin
                      state <= 3'h2;
                    end
                  end
                end
              end
            end
          end else begin
            if(T_145) begin
              if(T_203) begin
                if(isHi) begin
                  state <= 3'h3;
                end else begin
                  state <= 3'h5;
                end
              end else begin
                if(T_141) begin
                  if(neg_out) begin
                    state <= 3'h4;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_140) begin
                    state <= 3'h5;
                  end else begin
                    if(T_135) begin
                      state <= 3'h2;
                    end
                  end
                end
              end
            end else begin
              if(T_141) begin
                state <= T_143;
              end else begin
                if(T_140) begin
                  state <= 3'h5;
                end else begin
                  if(T_135) begin
                    state <= 3'h2;
                  end
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        req_fn <= io_req_bits_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        req_dw <= io_req_bits_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        req_in1 <= io_req_bits_in1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        req_in2 <= io_req_bits_in2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        count <= {{6'd0}, 1'h0};
      end else begin
        if(T_208) begin
          if(T_614) begin
            count <= {{1'd0}, T_619};
          end else begin
            count <= T_200;
          end
        end else begin
          if(T_145) begin
            count <= T_200;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        neg_out <= T_644;
      end else begin
        if(T_208) begin
          if(T_629) begin
            neg_out <= 1'h0;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        isMul <= T_71;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        isHi <= T_83;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        divisor <= T_645;
      end else begin
        if(T_135) begin
          if(T_139) begin
            divisor <= subtractor;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_633) begin
        remainder <= {{66'd0}, lhs_in};
      end else begin
        if(T_208) begin
          remainder <= {{1'd0}, GEN_14};
        end else begin
          if(T_145) begin
            remainder <= T_197;
          end else begin
            if(T_141) begin
              remainder <= {{66'd0}, T_142};
            end else begin
              if(T_140) begin
                remainder <= {{66'd0}, negated_remainder};
              end else begin
                if(T_135) begin
                  if(T_137) begin
                    remainder <= {{66'd0}, negated_remainder};
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module Rocket(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip,
  output  io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output  io_imem_resp_ready,
  input   io_imem_resp_valid,
  input  [39:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data_0,
  input   io_imem_resp_bits_mask,
  input   io_imem_resp_bits_xcpt_if,
  input   io_imem_btb_resp_valid,
  input   io_imem_btb_resp_bits_taken,
  input   io_imem_btb_resp_bits_mask,
  input   io_imem_btb_resp_bits_bridx,
  input  [38:0] io_imem_btb_resp_bits_target,
  input  [5:0] io_imem_btb_resp_bits_entry,
  input  [6:0] io_imem_btb_resp_bits_bht_history,
  input  [1:0] io_imem_btb_resp_bits_bht_value,
  output  io_imem_btb_update_valid,
  output  io_imem_btb_update_bits_prediction_valid,
  output  io_imem_btb_update_bits_prediction_bits_taken,
  output  io_imem_btb_update_bits_prediction_bits_mask,
  output  io_imem_btb_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_btb_update_bits_prediction_bits_target,
  output [5:0] io_imem_btb_update_bits_prediction_bits_entry,
  output [6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
  output [38:0] io_imem_btb_update_bits_pc,
  output [38:0] io_imem_btb_update_bits_target,
  output  io_imem_btb_update_bits_taken,
  output  io_imem_btb_update_bits_isJump,
  output  io_imem_btb_update_bits_isReturn,
  output [38:0] io_imem_btb_update_bits_br_pc,
  output  io_imem_bht_update_valid,
  output  io_imem_bht_update_bits_prediction_valid,
  output  io_imem_bht_update_bits_prediction_bits_taken,
  output  io_imem_bht_update_bits_prediction_bits_mask,
  output  io_imem_bht_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_bht_update_bits_prediction_bits_target,
  output [5:0] io_imem_bht_update_bits_prediction_bits_entry,
  output [6:0] io_imem_bht_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
  output [38:0] io_imem_bht_update_bits_pc,
  output  io_imem_bht_update_bits_taken,
  output  io_imem_bht_update_bits_mispredict,
  output  io_imem_ras_update_valid,
  output  io_imem_ras_update_bits_isCall,
  output  io_imem_ras_update_bits_isReturn,
  output [38:0] io_imem_ras_update_bits_returnAddr,
  output  io_imem_ras_update_bits_prediction_valid,
  output  io_imem_ras_update_bits_prediction_bits_taken,
  output  io_imem_ras_update_bits_prediction_bits_mask,
  output  io_imem_ras_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_ras_update_bits_prediction_bits_target,
  output [5:0] io_imem_ras_update_bits_prediction_bits_entry,
  output [6:0] io_imem_ras_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
  output  io_imem_flush_icache,
  output  io_imem_flush_tlb,
  input  [39:0] io_imem_npc,
  input   io_dmem_req_ready,
  output  io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [8:0] io_dmem_req_bits_tag,
  output [4:0] io_dmem_req_bits_cmd,
  output [2:0] io_dmem_req_bits_typ,
  output  io_dmem_req_bits_phys,
  output [63:0] io_dmem_req_bits_data,
  output  io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data,
  input   io_dmem_s2_nack,
  input   io_dmem_resp_valid,
  input  [39:0] io_dmem_resp_bits_addr,
  input  [8:0] io_dmem_resp_bits_tag,
  input  [4:0] io_dmem_resp_bits_cmd,
  input  [2:0] io_dmem_resp_bits_typ,
  input  [63:0] io_dmem_resp_bits_data,
  input   io_dmem_resp_bits_replay,
  input   io_dmem_resp_bits_has_data,
  input  [63:0] io_dmem_resp_bits_data_word_bypass,
  input  [63:0] io_dmem_resp_bits_store_data,
  input   io_dmem_replay_next,
  input   io_dmem_xcpt_ma_ld,
  input   io_dmem_xcpt_ma_st,
  input   io_dmem_xcpt_pf_ld,
  input   io_dmem_xcpt_pf_st,
  output  io_dmem_invalidate_lr,
  input   io_dmem_ordered,
  output [6:0] io_ptw_ptbr_asid,
  output [37:0] io_ptw_ptbr_ppn,
  output  io_ptw_invalidate,
  output  io_ptw_status_debug,
  output [1:0] io_ptw_status_prv,
  output  io_ptw_status_sd,
  output [30:0] io_ptw_status_zero3,
  output  io_ptw_status_sd_rv32,
  output [1:0] io_ptw_status_zero2,
  output [4:0] io_ptw_status_vm,
  output [4:0] io_ptw_status_zero1,
  output  io_ptw_status_pum,
  output  io_ptw_status_mprv,
  output [1:0] io_ptw_status_xs,
  output [1:0] io_ptw_status_fs,
  output [1:0] io_ptw_status_mpp,
  output [1:0] io_ptw_status_hpp,
  output  io_ptw_status_spp,
  output  io_ptw_status_mpie,
  output  io_ptw_status_hpie,
  output  io_ptw_status_spie,
  output  io_ptw_status_upie,
  output  io_ptw_status_mie,
  output  io_ptw_status_hie,
  output  io_ptw_status_sie,
  output  io_ptw_status_uie,
  output [31:0] io_fpu_inst,
  output [63:0] io_fpu_fromint_data,
  output [2:0] io_fpu_fcsr_rm,
  input   io_fpu_fcsr_flags_valid,
  input  [4:0] io_fpu_fcsr_flags_bits,
  input  [63:0] io_fpu_store_data,
  input  [63:0] io_fpu_toint_data,
  output  io_fpu_dmem_resp_val,
  output [2:0] io_fpu_dmem_resp_type,
  output [4:0] io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output  io_fpu_valid,
  input   io_fpu_fcsr_rdy,
  input   io_fpu_nack_mem,
  input   io_fpu_illegal_rm,
  output  io_fpu_killx,
  output  io_fpu_killm,
  input  [4:0] io_fpu_dec_cmd,
  input   io_fpu_dec_ldst,
  input   io_fpu_dec_wen,
  input   io_fpu_dec_ren1,
  input   io_fpu_dec_ren2,
  input   io_fpu_dec_ren3,
  input   io_fpu_dec_swap12,
  input   io_fpu_dec_swap23,
  input   io_fpu_dec_single,
  input   io_fpu_dec_fromint,
  input   io_fpu_dec_toint,
  input   io_fpu_dec_fastpipe,
  input   io_fpu_dec_fma,
  input   io_fpu_dec_div,
  input   io_fpu_dec_sqrt,
  input   io_fpu_dec_round,
  input   io_fpu_dec_wflags,
  input   io_fpu_sboard_set,
  input   io_fpu_sboard_clr,
  input  [4:0] io_fpu_sboard_clra,
  input   io_fpu_cp_req_ready,
  output  io_fpu_cp_req_valid,
  output [4:0] io_fpu_cp_req_bits_cmd,
  output  io_fpu_cp_req_bits_ldst,
  output  io_fpu_cp_req_bits_wen,
  output  io_fpu_cp_req_bits_ren1,
  output  io_fpu_cp_req_bits_ren2,
  output  io_fpu_cp_req_bits_ren3,
  output  io_fpu_cp_req_bits_swap12,
  output  io_fpu_cp_req_bits_swap23,
  output  io_fpu_cp_req_bits_single,
  output  io_fpu_cp_req_bits_fromint,
  output  io_fpu_cp_req_bits_toint,
  output  io_fpu_cp_req_bits_fastpipe,
  output  io_fpu_cp_req_bits_fma,
  output  io_fpu_cp_req_bits_div,
  output  io_fpu_cp_req_bits_sqrt,
  output  io_fpu_cp_req_bits_round,
  output  io_fpu_cp_req_bits_wflags,
  output [2:0] io_fpu_cp_req_bits_rm,
  output [1:0] io_fpu_cp_req_bits_typ,
  output [64:0] io_fpu_cp_req_bits_in1,
  output [64:0] io_fpu_cp_req_bits_in2,
  output [64:0] io_fpu_cp_req_bits_in3,
  output  io_fpu_cp_resp_ready,
  input   io_fpu_cp_resp_valid,
  input  [64:0] io_fpu_cp_resp_bits_data,
  input  [4:0] io_fpu_cp_resp_bits_exc,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [63:0] io_rocc_cmd_bits_rs1,
  output [63:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [63:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [39:0] io_rocc_mem_req_bits_addr,
  input  [8:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [63:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [63:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [39:0] io_rocc_mem_resp_bits_addr,
  output [8:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [63:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [63:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  output  io_rocc_status_debug,
  output [1:0] io_rocc_status_prv,
  output  io_rocc_status_sd,
  output [30:0] io_rocc_status_zero3,
  output  io_rocc_status_sd_rv32,
  output [1:0] io_rocc_status_zero2,
  output [4:0] io_rocc_status_vm,
  output [4:0] io_rocc_status_zero1,
  output  io_rocc_status_pum,
  output  io_rocc_status_mprv,
  output [1:0] io_rocc_status_xs,
  output [1:0] io_rocc_status_fs,
  output [1:0] io_rocc_status_mpp,
  output [1:0] io_rocc_status_hpp,
  output  io_rocc_status_spp,
  output  io_rocc_status_mpie,
  output  io_rocc_status_hpie,
  output  io_rocc_status_spie,
  output  io_rocc_status_upie,
  output  io_rocc_status_mie,
  output  io_rocc_status_hie,
  output  io_rocc_status_sie,
  output  io_rocc_status_uie,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input  [1:0] io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [11:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output [1:0] io_rocc_autl_grant_bits_client_xact_id,
  output [2:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception,
  output [11:0] io_rocc_csr_waddr,
  output [63:0] io_rocc_csr_wdata,
  output  io_rocc_csr_wen,
  output  io_rocc_host_id
);
  reg  ex_ctrl_legal;
  reg [31:0] GEN_290;
  reg  ex_ctrl_fp;
  reg [31:0] GEN_291;
  reg  ex_ctrl_rocc;
  reg [31:0] GEN_292;
  reg  ex_ctrl_branch;
  reg [31:0] GEN_293;
  reg  ex_ctrl_jal;
  reg [31:0] GEN_294;
  reg  ex_ctrl_jalr;
  reg [31:0] GEN_295;
  reg  ex_ctrl_rxs2;
  reg [31:0] GEN_296;
  reg  ex_ctrl_rxs1;
  reg [31:0] GEN_297;
  reg [1:0] ex_ctrl_sel_alu2;
  reg [31:0] GEN_298;
  reg [1:0] ex_ctrl_sel_alu1;
  reg [31:0] GEN_299;
  reg [2:0] ex_ctrl_sel_imm;
  reg [31:0] GEN_300;
  reg  ex_ctrl_alu_dw;
  reg [31:0] GEN_301;
  reg [3:0] ex_ctrl_alu_fn;
  reg [31:0] GEN_302;
  reg  ex_ctrl_mem;
  reg [31:0] GEN_303;
  reg [4:0] ex_ctrl_mem_cmd;
  reg [31:0] GEN_304;
  reg [2:0] ex_ctrl_mem_type;
  reg [31:0] GEN_305;
  reg  ex_ctrl_rfs1;
  reg [31:0] GEN_306;
  reg  ex_ctrl_rfs2;
  reg [31:0] GEN_307;
  reg  ex_ctrl_rfs3;
  reg [31:0] GEN_308;
  reg  ex_ctrl_wfd;
  reg [31:0] GEN_309;
  reg  ex_ctrl_div;
  reg [31:0] GEN_310;
  reg  ex_ctrl_wxd;
  reg [31:0] GEN_311;
  reg [2:0] ex_ctrl_csr;
  reg [31:0] GEN_312;
  reg  ex_ctrl_fence_i;
  reg [31:0] GEN_313;
  reg  ex_ctrl_fence;
  reg [31:0] GEN_314;
  reg  ex_ctrl_amo;
  reg [31:0] GEN_315;
  reg  mem_ctrl_legal;
  reg [31:0] GEN_316;
  reg  mem_ctrl_fp;
  reg [31:0] GEN_317;
  reg  mem_ctrl_rocc;
  reg [31:0] GEN_318;
  reg  mem_ctrl_branch;
  reg [31:0] GEN_319;
  reg  mem_ctrl_jal;
  reg [31:0] GEN_320;
  reg  mem_ctrl_jalr;
  reg [31:0] GEN_321;
  reg  mem_ctrl_rxs2;
  reg [31:0] GEN_322;
  reg  mem_ctrl_rxs1;
  reg [31:0] GEN_323;
  reg [1:0] mem_ctrl_sel_alu2;
  reg [31:0] GEN_324;
  reg [1:0] mem_ctrl_sel_alu1;
  reg [31:0] GEN_325;
  reg [2:0] mem_ctrl_sel_imm;
  reg [31:0] GEN_326;
  reg  mem_ctrl_alu_dw;
  reg [31:0] GEN_327;
  reg [3:0] mem_ctrl_alu_fn;
  reg [31:0] GEN_328;
  reg  mem_ctrl_mem;
  reg [31:0] GEN_329;
  reg [4:0] mem_ctrl_mem_cmd;
  reg [31:0] GEN_330;
  reg [2:0] mem_ctrl_mem_type;
  reg [31:0] GEN_331;
  reg  mem_ctrl_rfs1;
  reg [31:0] GEN_332;
  reg  mem_ctrl_rfs2;
  reg [31:0] GEN_333;
  reg  mem_ctrl_rfs3;
  reg [31:0] GEN_334;
  reg  mem_ctrl_wfd;
  reg [31:0] GEN_335;
  reg  mem_ctrl_div;
  reg [31:0] GEN_336;
  reg  mem_ctrl_wxd;
  reg [31:0] GEN_337;
  reg [2:0] mem_ctrl_csr;
  reg [31:0] GEN_338;
  reg  mem_ctrl_fence_i;
  reg [31:0] GEN_339;
  reg  mem_ctrl_fence;
  reg [31:0] GEN_340;
  reg  mem_ctrl_amo;
  reg [31:0] GEN_341;
  reg  wb_ctrl_legal;
  reg [31:0] GEN_342;
  reg  wb_ctrl_fp;
  reg [31:0] GEN_343;
  reg  wb_ctrl_rocc;
  reg [31:0] GEN_344;
  reg  wb_ctrl_branch;
  reg [31:0] GEN_345;
  reg  wb_ctrl_jal;
  reg [31:0] GEN_346;
  reg  wb_ctrl_jalr;
  reg [31:0] GEN_347;
  reg  wb_ctrl_rxs2;
  reg [31:0] GEN_348;
  reg  wb_ctrl_rxs1;
  reg [31:0] GEN_349;
  reg [1:0] wb_ctrl_sel_alu2;
  reg [31:0] GEN_350;
  reg [1:0] wb_ctrl_sel_alu1;
  reg [31:0] GEN_351;
  reg [2:0] wb_ctrl_sel_imm;
  reg [31:0] GEN_352;
  reg  wb_ctrl_alu_dw;
  reg [31:0] GEN_353;
  reg [3:0] wb_ctrl_alu_fn;
  reg [31:0] GEN_354;
  reg  wb_ctrl_mem;
  reg [31:0] GEN_355;
  reg [4:0] wb_ctrl_mem_cmd;
  reg [31:0] GEN_356;
  reg [2:0] wb_ctrl_mem_type;
  reg [31:0] GEN_357;
  reg  wb_ctrl_rfs1;
  reg [31:0] GEN_358;
  reg  wb_ctrl_rfs2;
  reg [31:0] GEN_359;
  reg  wb_ctrl_rfs3;
  reg [31:0] GEN_360;
  reg  wb_ctrl_wfd;
  reg [31:0] GEN_361;
  reg  wb_ctrl_div;
  reg [31:0] GEN_362;
  reg  wb_ctrl_wxd;
  reg [31:0] GEN_363;
  reg [2:0] wb_ctrl_csr;
  reg [31:0] GEN_364;
  reg  wb_ctrl_fence_i;
  reg [31:0] GEN_365;
  reg  wb_ctrl_fence;
  reg [31:0] GEN_366;
  reg  wb_ctrl_amo;
  reg [31:0] GEN_367;
  reg  ex_reg_xcpt_interrupt;
  reg [31:0] GEN_368;
  reg  ex_reg_valid;
  reg [31:0] GEN_369;
  reg  ex_reg_btb_hit;
  reg [31:0] GEN_370;
  reg  ex_reg_btb_resp_taken;
  reg [31:0] GEN_371;
  reg  ex_reg_btb_resp_mask;
  reg [31:0] GEN_372;
  reg  ex_reg_btb_resp_bridx;
  reg [31:0] GEN_373;
  reg [38:0] ex_reg_btb_resp_target;
  reg [63:0] GEN_374;
  reg [5:0] ex_reg_btb_resp_entry;
  reg [31:0] GEN_375;
  reg [6:0] ex_reg_btb_resp_bht_history;
  reg [31:0] GEN_376;
  reg [1:0] ex_reg_btb_resp_bht_value;
  reg [31:0] GEN_377;
  reg  ex_reg_xcpt;
  reg [31:0] GEN_378;
  reg  ex_reg_flush_pipe;
  reg [31:0] GEN_379;
  reg  ex_reg_load_use;
  reg [31:0] GEN_380;
  reg [63:0] ex_reg_cause;
  reg [63:0] GEN_381;
  reg [39:0] ex_reg_pc;
  reg [63:0] GEN_382;
  reg [31:0] ex_reg_inst;
  reg [31:0] GEN_383;
  reg  mem_reg_xcpt_interrupt;
  reg [31:0] GEN_384;
  reg  mem_reg_valid;
  reg [31:0] GEN_385;
  reg  mem_reg_btb_hit;
  reg [31:0] GEN_386;
  reg  mem_reg_btb_resp_taken;
  reg [31:0] GEN_387;
  reg  mem_reg_btb_resp_mask;
  reg [31:0] GEN_388;
  reg  mem_reg_btb_resp_bridx;
  reg [31:0] GEN_389;
  reg [38:0] mem_reg_btb_resp_target;
  reg [63:0] GEN_390;
  reg [5:0] mem_reg_btb_resp_entry;
  reg [31:0] GEN_391;
  reg [6:0] mem_reg_btb_resp_bht_history;
  reg [31:0] GEN_392;
  reg [1:0] mem_reg_btb_resp_bht_value;
  reg [31:0] GEN_393;
  reg  mem_reg_xcpt;
  reg [31:0] GEN_394;
  reg  mem_reg_replay;
  reg [31:0] GEN_395;
  reg  mem_reg_flush_pipe;
  reg [31:0] GEN_396;
  reg [63:0] mem_reg_cause;
  reg [63:0] GEN_397;
  reg  mem_reg_slow_bypass;
  reg [31:0] GEN_398;
  reg  mem_reg_load;
  reg [31:0] GEN_399;
  reg  mem_reg_store;
  reg [31:0] GEN_400;
  reg [39:0] mem_reg_pc;
  reg [63:0] GEN_401;
  reg [31:0] mem_reg_inst;
  reg [31:0] GEN_402;
  reg [63:0] mem_reg_wdata;
  reg [63:0] GEN_403;
  reg [63:0] mem_reg_rs2;
  reg [63:0] GEN_404;
  wire  take_pc_mem;
  reg  wb_reg_valid;
  reg [31:0] GEN_405;
  reg  wb_reg_xcpt;
  reg [31:0] GEN_406;
  reg  wb_reg_mem_xcpt;
  reg [31:0] GEN_407;
  reg  wb_reg_replay;
  reg [31:0] GEN_408;
  reg [63:0] wb_reg_cause;
  reg [63:0] GEN_409;
  reg [39:0] wb_reg_pc;
  reg [63:0] GEN_410;
  reg [31:0] wb_reg_inst;
  reg [31:0] GEN_411;
  reg [63:0] wb_reg_wdata;
  reg [63:0] GEN_412;
  reg [63:0] wb_reg_rs2;
  reg [63:0] GEN_413;
  wire  take_pc_wb;
  wire  take_pc_mem_wb;
  wire  id_ctrl_legal;
  wire  id_ctrl_fp;
  wire  id_ctrl_rocc;
  wire  id_ctrl_branch;
  wire  id_ctrl_jal;
  wire  id_ctrl_jalr;
  wire  id_ctrl_rxs2;
  wire  id_ctrl_rxs1;
  wire [1:0] id_ctrl_sel_alu2;
  wire [1:0] id_ctrl_sel_alu1;
  wire [2:0] id_ctrl_sel_imm;
  wire  id_ctrl_alu_dw;
  wire [3:0] id_ctrl_alu_fn;
  wire  id_ctrl_mem;
  wire [4:0] id_ctrl_mem_cmd;
  wire [2:0] id_ctrl_mem_type;
  wire  id_ctrl_rfs1;
  wire  id_ctrl_rfs2;
  wire  id_ctrl_rfs3;
  wire  id_ctrl_wfd;
  wire  id_ctrl_div;
  wire  id_ctrl_wxd;
  wire [2:0] id_ctrl_csr;
  wire  id_ctrl_fence_i;
  wire  id_ctrl_fence;
  wire  id_ctrl_amo;
  wire [31:0] T_6629;
  wire  T_6631;
  wire [31:0] T_6633;
  wire  T_6635;
  wire [31:0] T_6637;
  wire  T_6639;
  wire [31:0] T_6641;
  wire  T_6643;
  wire [31:0] T_6645;
  wire  T_6647;
  wire [31:0] T_6649;
  wire  T_6651;
  wire [31:0] T_6653;
  wire  T_6655;
  wire [31:0] T_6657;
  wire  T_6659;
  wire [31:0] T_6661;
  wire  T_6663;
  wire [31:0] T_6665;
  wire  T_6667;
  wire [31:0] T_6669;
  wire  T_6671;
  wire [31:0] T_6673;
  wire  T_6675;
  wire [31:0] T_6677;
  wire  T_6679;
  wire  T_6683;
  wire [31:0] T_6685;
  wire  T_6687;
  wire  T_6691;
  wire [31:0] T_6693;
  wire  T_6695;
  wire [31:0] T_6697;
  wire  T_6699;
  wire  T_6703;
  wire [31:0] T_6705;
  wire  T_6707;
  wire [31:0] T_6709;
  wire  T_6711;
  wire [31:0] T_6713;
  wire  T_6715;
  wire [31:0] T_6717;
  wire  T_6719;
  wire [31:0] T_6721;
  wire  T_6723;
  wire  T_6725;
  wire  T_6727;
  wire [31:0] T_6729;
  wire  T_6731;
  wire [31:0] T_6733;
  wire  T_6735;
  wire [31:0] T_6737;
  wire  T_6739;
  wire  T_6742;
  wire  T_6743;
  wire  T_6744;
  wire  T_6745;
  wire  T_6746;
  wire  T_6747;
  wire  T_6748;
  wire  T_6749;
  wire  T_6750;
  wire  T_6751;
  wire  T_6752;
  wire  T_6753;
  wire  T_6754;
  wire  T_6755;
  wire  T_6756;
  wire  T_6757;
  wire  T_6758;
  wire  T_6759;
  wire  T_6760;
  wire  T_6761;
  wire  T_6762;
  wire  T_6763;
  wire  T_6764;
  wire  T_6765;
  wire  T_6766;
  wire  T_6767;
  wire  T_6768;
  wire  T_6769;
  wire [31:0] T_6773;
  wire  T_6775;
  wire [31:0] T_6779;
  wire  T_6781;
  wire [31:0] T_6785;
  wire  T_6787;
  wire [31:0] T_6791;
  wire  T_6793;
  wire [31:0] T_6795;
  wire  T_6797;
  wire [31:0] T_6799;
  wire  T_6801;
  wire  T_6804;
  wire  T_6805;
  wire [31:0] T_6807;
  wire  T_6809;
  wire [31:0] T_6811;
  wire  T_6813;
  wire [31:0] T_6815;
  wire  T_6817;
  wire [31:0] T_6819;
  wire  T_6821;
  wire  T_6824;
  wire  T_6825;
  wire  T_6826;
  wire [31:0] T_6828;
  wire  T_6830;
  wire [31:0] T_6832;
  wire  T_6834;
  wire [31:0] T_6836;
  wire  T_6838;
  wire [31:0] T_6840;
  wire  T_6842;
  wire  T_6845;
  wire  T_6846;
  wire  T_6847;
  wire  T_6848;
  wire  T_6852;
  wire [31:0] T_6854;
  wire  T_6856;
  wire  T_6859;
  wire  T_6860;
  wire  T_6861;
  wire [1:0] T_6862;
  wire [31:0] T_6864;
  wire  T_6866;
  wire  T_6869;
  wire  T_6870;
  wire  T_6871;
  wire [31:0] T_6873;
  wire  T_6875;
  wire  T_6878;
  wire [1:0] T_6879;
  wire  T_6883;
  wire  T_6887;
  wire  T_6890;
  wire  T_6894;
  wire  T_6897;
  wire  T_6901;
  wire [31:0] T_6903;
  wire  T_6905;
  wire  T_6908;
  wire  T_6909;
  wire [1:0] T_6910;
  wire [2:0] T_6911;
  wire [31:0] T_6913;
  wire  T_6915;
  wire [31:0] T_6917;
  wire  T_6919;
  wire  T_6922;
  wire [31:0] T_6924;
  wire  T_6926;
  wire [31:0] T_6928;
  wire  T_6930;
  wire [31:0] T_6932;
  wire  T_6934;
  wire  T_6937;
  wire  T_6938;
  wire [31:0] T_6940;
  wire  T_6942;
  wire [31:0] T_6944;
  wire  T_6946;
  wire  T_6950;
  wire [31:0] T_6952;
  wire  T_6954;
  wire [31:0] T_6956;
  wire  T_6958;
  wire [31:0] T_6960;
  wire  T_6962;
  wire  T_6965;
  wire  T_6966;
  wire  T_6967;
  wire  T_6968;
  wire  T_6969;
  wire [31:0] T_6971;
  wire  T_6973;
  wire [31:0] T_6975;
  wire  T_6977;
  wire [31:0] T_6979;
  wire  T_6981;
  wire [31:0] T_6983;
  wire  T_6985;
  wire  T_6988;
  wire  T_6989;
  wire  T_6990;
  wire  T_6994;
  wire [31:0] T_6996;
  wire  T_6998;
  wire  T_7001;
  wire  T_7002;
  wire  T_7003;
  wire [1:0] T_7004;
  wire [2:0] T_7005;
  wire [3:0] T_7006;
  wire [31:0] T_7008;
  wire  T_7010;
  wire [31:0] T_7012;
  wire  T_7014;
  wire  T_7018;
  wire  T_7019;
  wire  T_7020;
  wire  T_7021;
  wire  T_7022;
  wire [31:0] T_7024;
  wire  T_7026;
  wire [31:0] T_7028;
  wire  T_7030;
  wire [31:0] T_7032;
  wire  T_7034;
  wire [31:0] T_7036;
  wire  T_7038;
  wire  T_7041;
  wire  T_7042;
  wire  T_7043;
  wire [31:0] T_7045;
  wire  T_7047;
  wire [31:0] T_7049;
  wire  T_7051;
  wire  T_7054;
  wire [31:0] T_7056;
  wire  T_7058;
  wire [31:0] T_7060;
  wire  T_7062;
  wire [31:0] T_7064;
  wire  T_7066;
  wire  T_7069;
  wire  T_7070;
  wire  T_7071;
  wire [31:0] T_7073;
  wire  T_7075;
  wire [1:0] T_7079;
  wire [2:0] T_7080;
  wire [3:0] T_7081;
  wire [4:0] T_7082;
  wire [31:0] T_7084;
  wire  T_7086;
  wire [31:0] T_7090;
  wire  T_7092;
  wire [31:0] T_7096;
  wire  T_7098;
  wire [1:0] T_7101;
  wire [2:0] T_7102;
  wire [31:0] T_7108;
  wire  T_7110;
  wire  T_7116;
  wire [31:0] T_7118;
  wire  T_7120;
  wire  T_7124;
  wire [31:0] T_7126;
  wire  T_7128;
  wire  T_7132;
  wire  T_7135;
  wire  T_7136;
  wire  T_7137;
  wire  T_7138;
  wire  T_7139;
  wire  T_7140;
  wire [31:0] T_7142;
  wire  T_7144;
  wire  T_7150;
  wire [31:0] T_7154;
  wire  T_7156;
  wire [1:0] T_7159;
  wire [2:0] T_7160;
  wire [31:0] T_7162;
  wire  T_7164;
  wire  T_7170;
  wire [31:0] T_7174;
  wire  T_7176;
  wire [4:0] id_raddr3;
  wire [4:0] id_raddr2;
  wire [4:0] id_raddr1;
  wire [4:0] id_waddr;
  wire  id_load_use;
  reg  id_reg_fence;
  reg [31:0] GEN_414;
  reg [63:0] T_7183 [0:30];
  reg [63:0] GEN_415;
  wire [63:0] T_7183_T_7193_data;
  wire [4:0] T_7183_T_7193_addr;
  wire  T_7183_T_7193_en;
  wire [63:0] T_7183_T_7204_data;
  wire [4:0] T_7183_T_7204_addr;
  wire  T_7183_T_7204_en;
  wire [63:0] T_7183_T_7850_data;
  wire [4:0] T_7183_T_7850_addr;
  wire  T_7183_T_7850_mask;
  wire  T_7183_T_7850_en;
  wire [63:0] T_7185;
  wire [4:0] GEN_170;
  wire  T_7188;
  wire [4:0] T_7192;
  wire [63:0] T_7194;
  wire [63:0] T_7196;
  wire [4:0] T_7203;
  wire [63:0] T_7205;
  wire  ctrl_killd;
  wire  csr_clk;
  wire  csr_reset;
  wire  csr_io_prci_reset;
  wire  csr_io_prci_id;
  wire  csr_io_prci_interrupts_meip;
  wire  csr_io_prci_interrupts_seip;
  wire  csr_io_prci_interrupts_debug;
  wire  csr_io_prci_interrupts_mtip;
  wire  csr_io_prci_interrupts_msip;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [63:0] csr_io_rw_rdata;
  wire [63:0] csr_io_rw_wdata;
  wire  csr_io_csr_stall;
  wire  csr_io_csr_xcpt;
  wire  csr_io_eret;
  wire  csr_io_singleStep;
  wire  csr_io_status_debug;
  wire [1:0] csr_io_status_prv;
  wire  csr_io_status_sd;
  wire [30:0] csr_io_status_zero3;
  wire  csr_io_status_sd_rv32;
  wire [1:0] csr_io_status_zero2;
  wire [4:0] csr_io_status_vm;
  wire [4:0] csr_io_status_zero1;
  wire  csr_io_status_pum;
  wire  csr_io_status_mprv;
  wire [1:0] csr_io_status_xs;
  wire [1:0] csr_io_status_fs;
  wire [1:0] csr_io_status_mpp;
  wire [1:0] csr_io_status_hpp;
  wire  csr_io_status_spp;
  wire  csr_io_status_mpie;
  wire  csr_io_status_hpie;
  wire  csr_io_status_spie;
  wire  csr_io_status_upie;
  wire  csr_io_status_mie;
  wire  csr_io_status_hie;
  wire  csr_io_status_sie;
  wire  csr_io_status_uie;
  wire [6:0] csr_io_ptbr_asid;
  wire [37:0] csr_io_ptbr_ppn;
  wire [39:0] csr_io_evec;
  wire  csr_io_exception;
  wire  csr_io_retire;
  wire  csr_io_uarch_counters_0;
  wire  csr_io_uarch_counters_1;
  wire  csr_io_uarch_counters_2;
  wire  csr_io_uarch_counters_3;
  wire  csr_io_uarch_counters_4;
  wire  csr_io_uarch_counters_5;
  wire  csr_io_uarch_counters_6;
  wire  csr_io_uarch_counters_7;
  wire  csr_io_uarch_counters_8;
  wire  csr_io_uarch_counters_9;
  wire  csr_io_uarch_counters_10;
  wire  csr_io_uarch_counters_11;
  wire  csr_io_uarch_counters_12;
  wire  csr_io_uarch_counters_13;
  wire  csr_io_uarch_counters_14;
  wire  csr_io_uarch_counters_15;
  wire [63:0] csr_io_cause;
  wire [39:0] csr_io_pc;
  wire [39:0] csr_io_badaddr;
  wire  csr_io_fatc;
  wire [63:0] csr_io_time;
  wire [2:0] csr_io_fcsr_rm;
  wire  csr_io_fcsr_flags_valid;
  wire [4:0] csr_io_fcsr_flags_bits;
  wire  csr_io_rocc_cmd_ready;
  wire  csr_io_rocc_cmd_valid;
  wire [6:0] csr_io_rocc_cmd_bits_inst_funct;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs1;
  wire  csr_io_rocc_cmd_bits_inst_xd;
  wire  csr_io_rocc_cmd_bits_inst_xs1;
  wire  csr_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rd;
  wire [6:0] csr_io_rocc_cmd_bits_inst_opcode;
  wire [63:0] csr_io_rocc_cmd_bits_rs1;
  wire [63:0] csr_io_rocc_cmd_bits_rs2;
  wire  csr_io_rocc_resp_ready;
  wire  csr_io_rocc_resp_valid;
  wire [4:0] csr_io_rocc_resp_bits_rd;
  wire [63:0] csr_io_rocc_resp_bits_data;
  wire  csr_io_rocc_mem_req_ready;
  wire  csr_io_rocc_mem_req_valid;
  wire [39:0] csr_io_rocc_mem_req_bits_addr;
  wire [8:0] csr_io_rocc_mem_req_bits_tag;
  wire [4:0] csr_io_rocc_mem_req_bits_cmd;
  wire [2:0] csr_io_rocc_mem_req_bits_typ;
  wire  csr_io_rocc_mem_req_bits_phys;
  wire [63:0] csr_io_rocc_mem_req_bits_data;
  wire  csr_io_rocc_mem_s1_kill;
  wire [63:0] csr_io_rocc_mem_s1_data;
  wire  csr_io_rocc_mem_s2_nack;
  wire  csr_io_rocc_mem_resp_valid;
  wire [39:0] csr_io_rocc_mem_resp_bits_addr;
  wire [8:0] csr_io_rocc_mem_resp_bits_tag;
  wire [4:0] csr_io_rocc_mem_resp_bits_cmd;
  wire [2:0] csr_io_rocc_mem_resp_bits_typ;
  wire [63:0] csr_io_rocc_mem_resp_bits_data;
  wire  csr_io_rocc_mem_resp_bits_replay;
  wire  csr_io_rocc_mem_resp_bits_has_data;
  wire [63:0] csr_io_rocc_mem_resp_bits_data_word_bypass;
  wire [63:0] csr_io_rocc_mem_resp_bits_store_data;
  wire  csr_io_rocc_mem_replay_next;
  wire  csr_io_rocc_mem_xcpt_ma_ld;
  wire  csr_io_rocc_mem_xcpt_ma_st;
  wire  csr_io_rocc_mem_xcpt_pf_ld;
  wire  csr_io_rocc_mem_xcpt_pf_st;
  wire  csr_io_rocc_mem_invalidate_lr;
  wire  csr_io_rocc_mem_ordered;
  wire  csr_io_rocc_busy;
  wire  csr_io_rocc_status_debug;
  wire [1:0] csr_io_rocc_status_prv;
  wire  csr_io_rocc_status_sd;
  wire [30:0] csr_io_rocc_status_zero3;
  wire  csr_io_rocc_status_sd_rv32;
  wire [1:0] csr_io_rocc_status_zero2;
  wire [4:0] csr_io_rocc_status_vm;
  wire [4:0] csr_io_rocc_status_zero1;
  wire  csr_io_rocc_status_pum;
  wire  csr_io_rocc_status_mprv;
  wire [1:0] csr_io_rocc_status_xs;
  wire [1:0] csr_io_rocc_status_fs;
  wire [1:0] csr_io_rocc_status_mpp;
  wire [1:0] csr_io_rocc_status_hpp;
  wire  csr_io_rocc_status_spp;
  wire  csr_io_rocc_status_mpie;
  wire  csr_io_rocc_status_hpie;
  wire  csr_io_rocc_status_spie;
  wire  csr_io_rocc_status_upie;
  wire  csr_io_rocc_status_mie;
  wire  csr_io_rocc_status_hie;
  wire  csr_io_rocc_status_sie;
  wire  csr_io_rocc_status_uie;
  wire  csr_io_rocc_interrupt;
  wire  csr_io_rocc_autl_acquire_ready;
  wire  csr_io_rocc_autl_acquire_valid;
  wire [25:0] csr_io_rocc_autl_acquire_bits_addr_block;
  wire [1:0] csr_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] csr_io_rocc_autl_acquire_bits_addr_beat;
  wire  csr_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] csr_io_rocc_autl_acquire_bits_a_type;
  wire [11:0] csr_io_rocc_autl_acquire_bits_union;
  wire [63:0] csr_io_rocc_autl_acquire_bits_data;
  wire  csr_io_rocc_autl_grant_ready;
  wire  csr_io_rocc_autl_grant_valid;
  wire [2:0] csr_io_rocc_autl_grant_bits_addr_beat;
  wire [1:0] csr_io_rocc_autl_grant_bits_client_xact_id;
  wire [2:0] csr_io_rocc_autl_grant_bits_manager_xact_id;
  wire  csr_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] csr_io_rocc_autl_grant_bits_g_type;
  wire [63:0] csr_io_rocc_autl_grant_bits_data;
  wire  csr_io_rocc_fpu_req_ready;
  wire  csr_io_rocc_fpu_req_valid;
  wire [4:0] csr_io_rocc_fpu_req_bits_cmd;
  wire  csr_io_rocc_fpu_req_bits_ldst;
  wire  csr_io_rocc_fpu_req_bits_wen;
  wire  csr_io_rocc_fpu_req_bits_ren1;
  wire  csr_io_rocc_fpu_req_bits_ren2;
  wire  csr_io_rocc_fpu_req_bits_ren3;
  wire  csr_io_rocc_fpu_req_bits_swap12;
  wire  csr_io_rocc_fpu_req_bits_swap23;
  wire  csr_io_rocc_fpu_req_bits_single;
  wire  csr_io_rocc_fpu_req_bits_fromint;
  wire  csr_io_rocc_fpu_req_bits_toint;
  wire  csr_io_rocc_fpu_req_bits_fastpipe;
  wire  csr_io_rocc_fpu_req_bits_fma;
  wire  csr_io_rocc_fpu_req_bits_div;
  wire  csr_io_rocc_fpu_req_bits_sqrt;
  wire  csr_io_rocc_fpu_req_bits_round;
  wire  csr_io_rocc_fpu_req_bits_wflags;
  wire [2:0] csr_io_rocc_fpu_req_bits_rm;
  wire [1:0] csr_io_rocc_fpu_req_bits_typ;
  wire [64:0] csr_io_rocc_fpu_req_bits_in1;
  wire [64:0] csr_io_rocc_fpu_req_bits_in2;
  wire [64:0] csr_io_rocc_fpu_req_bits_in3;
  wire  csr_io_rocc_fpu_resp_ready;
  wire  csr_io_rocc_fpu_resp_valid;
  wire [64:0] csr_io_rocc_fpu_resp_bits_data;
  wire [4:0] csr_io_rocc_fpu_resp_bits_exc;
  wire  csr_io_rocc_exception;
  wire [11:0] csr_io_rocc_csr_waddr;
  wire [63:0] csr_io_rocc_csr_wdata;
  wire  csr_io_rocc_csr_wen;
  wire  csr_io_rocc_host_id;
  wire  csr_io_interrupt;
  wire [63:0] csr_io_interrupt_cause;
  wire [3:0] csr_io_bp_0_control_tdrtype;
  wire [4:0] csr_io_bp_0_control_bpamaskmax;
  wire [35:0] csr_io_bp_0_control_reserved;
  wire [7:0] csr_io_bp_0_control_bpaction;
  wire [3:0] csr_io_bp_0_control_bpmatch;
  wire  csr_io_bp_0_control_m;
  wire  csr_io_bp_0_control_h;
  wire  csr_io_bp_0_control_s;
  wire  csr_io_bp_0_control_u;
  wire  csr_io_bp_0_control_r;
  wire  csr_io_bp_0_control_w;
  wire  csr_io_bp_0_control_x;
  wire [38:0] csr_io_bp_0_address;
  wire  id_csr_en;
  wire  id_system_insn;
  wire  T_7207;
  wire  T_7208;
  wire  T_7209;
  wire  id_csr_ren;
  wire [2:0] id_csr;
  wire [11:0] id_csr_addr;
  wire  T_7213;
  wire  T_7214;
  wire [11:0] T_7268;
  wire  T_7270;
  wire [11:0] T_7272;
  wire  T_7274;
  wire  T_7277;
  wire  T_7280;
  wire  T_7281;
  wire  id_csr_flush;
  wire  T_7283;
  wire [1:0] GEN_173;
  wire  T_7285;
  wire  T_7287;
  wire  T_7288;
  wire  T_7289;
  wire  T_7291;
  wire  T_7293;
  wire  T_7294;
  wire  id_illegal_insn;
  wire  id_amo_aq;
  wire  id_amo_rl;
  wire  T_7295;
  wire  id_fence_next;
  wire  T_7297;
  wire  id_mem_busy;
  wire  T_7303;
  wire  T_7305;
  wire  T_7306;
  wire  T_7308;
  wire  T_7309;
  wire  T_7310;
  wire  T_7311;
  wire  T_7312;
  wire  T_7313;
  wire  T_7314;
  wire  bpu_clk;
  wire  bpu_reset;
  wire  bpu_io_status_debug;
  wire [1:0] bpu_io_status_prv;
  wire  bpu_io_status_sd;
  wire [30:0] bpu_io_status_zero3;
  wire  bpu_io_status_sd_rv32;
  wire [1:0] bpu_io_status_zero2;
  wire [4:0] bpu_io_status_vm;
  wire [4:0] bpu_io_status_zero1;
  wire  bpu_io_status_pum;
  wire  bpu_io_status_mprv;
  wire [1:0] bpu_io_status_xs;
  wire [1:0] bpu_io_status_fs;
  wire [1:0] bpu_io_status_mpp;
  wire [1:0] bpu_io_status_hpp;
  wire  bpu_io_status_spp;
  wire  bpu_io_status_mpie;
  wire  bpu_io_status_hpie;
  wire  bpu_io_status_spie;
  wire  bpu_io_status_upie;
  wire  bpu_io_status_mie;
  wire  bpu_io_status_hie;
  wire  bpu_io_status_sie;
  wire  bpu_io_status_uie;
  wire [3:0] bpu_io_bp_0_control_tdrtype;
  wire [4:0] bpu_io_bp_0_control_bpamaskmax;
  wire [35:0] bpu_io_bp_0_control_reserved;
  wire [7:0] bpu_io_bp_0_control_bpaction;
  wire [3:0] bpu_io_bp_0_control_bpmatch;
  wire  bpu_io_bp_0_control_m;
  wire  bpu_io_bp_0_control_h;
  wire  bpu_io_bp_0_control_s;
  wire  bpu_io_bp_0_control_u;
  wire  bpu_io_bp_0_control_r;
  wire  bpu_io_bp_0_control_w;
  wire  bpu_io_bp_0_control_x;
  wire [38:0] bpu_io_bp_0_address;
  wire [38:0] bpu_io_pc;
  wire [38:0] bpu_io_ea;
  wire  bpu_io_xcpt_if;
  wire  bpu_io_xcpt_ld;
  wire  bpu_io_xcpt_st;
  wire  T_7318;
  wire  T_7319;
  wire  id_xcpt;
  wire [1:0] T_7320;
  wire [1:0] T_7321;
  wire [63:0] id_cause;
  wire [4:0] ex_waddr;
  wire [4:0] mem_waddr;
  wire [4:0] wb_waddr;
  wire  T_7325;
  wire  T_7326;
  wire  T_7328;
  wire  T_7329;
  wire  T_7331;
  wire  T_7333;
  wire  T_7334;
  wire  T_7335;
  wire  T_7336;
  wire  T_7338;
  wire  T_7339;
  wire  T_7341;
  wire  T_7342;
  wire  T_7343;
  wire  T_7344;
  wire  T_7346;
  wire [63:0] bypass_mux_0;
  wire [63:0] bypass_mux_1;
  wire [63:0] bypass_mux_2;
  wire [63:0] bypass_mux_3;
  reg  ex_reg_rs_bypass_0;
  reg [31:0] GEN_416;
  reg  ex_reg_rs_bypass_1;
  reg [31:0] GEN_417;
  reg [1:0] ex_reg_rs_lsb_0;
  reg [31:0] GEN_418;
  reg [1:0] ex_reg_rs_lsb_1;
  reg [31:0] GEN_419;
  reg [61:0] ex_reg_rs_msb_0;
  reg [63:0] GEN_420;
  reg [61:0] ex_reg_rs_msb_1;
  reg [63:0] GEN_421;
  wire [63:0] T_7374;
  wire [63:0] GEN_0;
  wire [1:0] GEN_177;
  wire [63:0] GEN_2;
  wire [63:0] GEN_3;
  wire [63:0] GEN_4;
  wire [63:0] T_7375;
  wire [63:0] T_7376;
  wire [63:0] GEN_1;
  wire [63:0] GEN_5;
  wire [63:0] GEN_6;
  wire [63:0] GEN_7;
  wire [63:0] T_7377;
  wire  T_7378;
  wire  T_7380;
  wire  T_7381;
  wire  T_7382;
  wire  T_7383;
  wire [10:0] T_7384;
  wire [10:0] T_7385;
  wire [10:0] T_7386;
  wire  T_7387;
  wire  T_7388;
  wire  T_7389;
  wire [7:0] T_7390;
  wire [7:0] T_7391;
  wire [7:0] T_7392;
  wire  T_7395;
  wire  T_7397;
  wire  T_7398;
  wire  T_7399;
  wire  T_7400;
  wire  T_7401;
  wire  T_7402;
  wire  T_7403;
  wire  T_7404;
  wire  T_7405;
  wire [5:0] T_7410;
  wire [5:0] T_7411;
  wire  T_7414;
  wire  T_7416;
  wire [3:0] T_7417;
  wire [3:0] T_7419;
  wire [3:0] T_7420;
  wire [3:0] T_7421;
  wire [3:0] T_7422;
  wire [3:0] T_7423;
  wire  T_7426;
  wire  T_7429;
  wire  T_7432;
  wire  T_7434;
  wire  T_7436;
  wire [9:0] T_7437;
  wire [10:0] T_7438;
  wire  T_7439;
  wire [7:0] T_7440;
  wire [8:0] T_7441;
  wire [10:0] T_7442;
  wire  T_7443;
  wire [11:0] T_7444;
  wire [20:0] T_7445;
  wire [31:0] T_7446;
  wire [31:0] ex_imm;
  wire [63:0] T_7448;
  wire [39:0] T_7449;
  wire  T_7450;
  wire  GEN_179;
  wire [39:0] T_7451;
  wire  T_7452;
  wire [63:0] ex_op1;
  wire [63:0] T_7454;
  wire  T_7456;
  wire [3:0] T_7457;
  wire  T_7458;
  wire [31:0] T_7459;
  wire  T_7460;
  wire [63:0] ex_op2;
  wire  alu_clk;
  wire  alu_reset;
  wire  alu_io_dw;
  wire [3:0] alu_io_fn;
  wire [63:0] alu_io_in2;
  wire [63:0] alu_io_in1;
  wire [63:0] alu_io_out;
  wire [63:0] alu_io_adder_out;
  wire  alu_io_cmp_out;
  wire [63:0] T_7461;
  wire [63:0] T_7462;
  wire  div_clk;
  wire  div_reset;
  wire  div_io_req_ready;
  wire  div_io_req_valid;
  wire [3:0] div_io_req_bits_fn;
  wire  div_io_req_bits_dw;
  wire [63:0] div_io_req_bits_in1;
  wire [63:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire  div_io_kill;
  wire  div_io_resp_ready;
  wire  div_io_resp_valid;
  wire [63:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire  T_7463;
  wire  T_7465;
  wire  T_7468;
  wire  T_7470;
  wire  T_7471;
  wire  T_7472;
  wire [63:0] GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire [38:0] GEN_12;
  wire [5:0] GEN_13;
  wire [6:0] GEN_14;
  wire [1:0] GEN_15;
  wire  T_7475;
  wire  T_7476;
  wire  T_7477;
  wire  GEN_16;
  wire  GEN_17;
  wire  T_7480;
  wire  T_7481;
  wire  T_7482;
  wire [1:0] T_7487;
  wire [1:0] T_7488;
  wire [1:0] T_7489;
  wire  T_7491;
  wire  T_7492;
  wire [1:0] T_7493;
  wire [61:0] T_7494;
  wire [1:0] GEN_18;
  wire [61:0] GEN_19;
  wire  T_7495;
  wire  T_7496;
  wire  T_7497;
  wire [1:0] T_7502;
  wire [1:0] T_7503;
  wire [1:0] T_7504;
  wire  T_7506;
  wire  T_7507;
  wire [1:0] T_7508;
  wire [61:0] T_7509;
  wire [1:0] GEN_20;
  wire [61:0] GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire [1:0] GEN_30;
  wire [1:0] GEN_31;
  wire [2:0] GEN_32;
  wire  GEN_33;
  wire [3:0] GEN_34;
  wire  GEN_35;
  wire [4:0] GEN_36;
  wire [2:0] GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire [2:0] GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire [38:0] GEN_52;
  wire [5:0] GEN_53;
  wire [6:0] GEN_54;
  wire [1:0] GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire [1:0] GEN_59;
  wire [61:0] GEN_60;
  wire  GEN_61;
  wire [1:0] GEN_62;
  wire [61:0] GEN_63;
  wire  T_7512;
  wire [31:0] GEN_64;
  wire [39:0] GEN_65;
  wire  ex_pc_valid;
  wire  T_7514;
  wire  wb_dcache_miss;
  wire  T_7516;
  wire  T_7517;
  wire  T_7519;
  wire  T_7520;
  wire  replay_ex_structural;
  wire  replay_ex_load_use;
  wire  T_7521;
  wire  replay_ex;
  wire  T_7522;
  wire  T_7524;
  wire  ctrl_killx;
  wire  T_7525;
  wire [2:0] T_7531_0;
  wire [2:0] T_7531_1;
  wire [2:0] T_7531_2;
  wire [2:0] T_7531_3;
  wire  T_7533;
  wire  T_7534;
  wire  T_7535;
  wire  T_7536;
  wire  T_7539;
  wire  T_7540;
  wire  T_7541;
  wire  ex_slow_bypass;
  wire  T_7542;
  wire  T_7543;
  wire  ex_xcpt;
  wire [63:0] ex_cause;
  wire  mem_br_taken;
  wire [39:0] T_7545;
  wire  T_7546;
  wire  T_7549;
  wire  T_7550;
  wire  T_7551;
  wire [10:0] T_7553;
  wire [10:0] T_7554;
  wire [10:0] T_7555;
  wire [7:0] T_7559;
  wire [7:0] T_7560;
  wire [7:0] T_7561;
  wire  T_7567;
  wire  T_7568;
  wire  T_7570;
  wire  T_7571;
  wire  T_7572;
  wire  T_7573;
  wire  T_7574;
  wire [5:0] T_7579;
  wire [3:0] T_7586;
  wire [3:0] T_7589;
  wire [9:0] T_7606;
  wire [10:0] T_7607;
  wire  T_7608;
  wire [7:0] T_7609;
  wire [8:0] T_7610;
  wire [10:0] T_7611;
  wire  T_7612;
  wire [11:0] T_7613;
  wire [20:0] T_7614;
  wire [31:0] T_7615;
  wire [31:0] T_7616;
  wire [7:0] T_7631;
  wire  T_7642;
  wire  T_7643;
  wire  T_7644;
  wire [9:0] T_7676;
  wire [10:0] T_7677;
  wire  T_7678;
  wire [7:0] T_7679;
  wire [8:0] T_7680;
  wire [20:0] T_7684;
  wire [31:0] T_7685;
  wire [31:0] T_7686;
  wire [3:0] GEN_181;
  wire [31:0] T_7688;
  wire [31:0] T_7689;
  wire [39:0] GEN_182;
  wire [40:0] T_7690;
  wire [39:0] T_7691;
  wire [39:0] mem_br_target;
  wire [63:0] T_7692;
  wire [63:0] T_7693;
  wire [63:0] mem_int_wdata;
  wire [25:0] T_7694;
  wire [1:0] T_7695;
  wire [1:0] T_7696;
  wire [25:0] GEN_183;
  wire  T_7698;
  wire [25:0] GEN_184;
  wire  T_7700;
  wire  T_7701;
  wire [1:0] GEN_186;
  wire  T_7703;
  wire [25:0] T_7704;
  wire  GEN_187;
  wire [25:0] GEN_188;
  wire  T_7706;
  wire [1:0] GEN_189;
  wire [25:0] GEN_190;
  wire  T_7709;
  wire  T_7710;
  wire [1:0] GEN_192;
  wire  T_7712;
  wire  T_7713;
  wire  T_7714;
  wire  T_7715;
  wire [38:0] T_7716;
  wire [39:0] T_7717;
  wire [39:0] T_7718;
  wire [39:0] T_7719;
  wire [39:0] GEN_194;
  wire [39:0] T_7721;
  wire [39:0] T_7722;
  wire [39:0] mem_npc;
  wire  T_7723;
  wire  T_7724;
  wire  T_7726;
  wire  mem_wrong_npc;
  wire  mem_npc_misaligned;
  wire  T_7729;
  wire  mem_cfi_taken;
  wire  T_7730;
  wire  want_take_pc_mem;
  wire  T_7732;
  wire  T_7733;
  wire  T_7735;
  wire  T_7738;
  wire  T_7741;
  wire  T_7744;
  wire [63:0] GEN_66;
  wire  T_7745;
  wire  T_7746;
  wire  T_7747;
  wire  T_7749;
  wire  T_7750;
  wire  T_7751;
  wire  T_7752;
  wire  T_7753;
  wire  T_7754;
  wire  T_7755;
  wire  T_7757;
  wire  T_7761;
  wire  T_7762;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire [38:0] GEN_70;
  wire [5:0] GEN_71;
  wire [6:0] GEN_72;
  wire [1:0] GEN_73;
  wire  T_7763;
  wire  T_7764;
  wire [63:0] GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire [1:0] GEN_83;
  wire [1:0] GEN_84;
  wire [2:0] GEN_85;
  wire  GEN_86;
  wire [3:0] GEN_87;
  wire  GEN_88;
  wire [4:0] GEN_89;
  wire [2:0] GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire [38:0] GEN_107;
  wire [5:0] GEN_108;
  wire [6:0] GEN_109;
  wire [1:0] GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire [31:0] GEN_113;
  wire [39:0] GEN_114;
  wire [63:0] GEN_115;
  wire [63:0] GEN_116;
  wire  T_7765;
  wire  T_7767;
  wire  T_7769;
  wire  T_7771;
  wire  T_7773;
  wire  T_7775;
  wire  T_7777;
  wire  T_7779;
  wire  T_7780;
  wire  T_7781;
  wire  T_7782;
  wire  T_7783;
  wire  mem_new_xcpt;
  wire [2:0] T_7784;
  wire [2:0] T_7785;
  wire [2:0] T_7786;
  wire [2:0] T_7787;
  wire [2:0] T_7788;
  wire [2:0] mem_new_cause;
  wire  T_7789;
  wire  T_7790;
  wire  mem_xcpt;
  wire [63:0] mem_cause;
  wire  dcache_kill_mem;
  wire  T_7792;
  wire  fpu_kill_mem;
  wire  T_7793;
  wire  replay_mem;
  wire  T_7794;
  wire  T_7795;
  wire  T_7797;
  wire  killm_common;
  wire  T_7798;
  reg  T_7799;
  reg [31:0] GEN_422;
  wire  T_7800;
  wire  T_7801;
  wire  ctrl_killm;
  wire  T_7803;
  wire  T_7805;
  wire  T_7806;
  wire  T_7809;
  wire  T_7813;
  wire  T_7814;
  wire [63:0] GEN_117;
  wire  T_7815;
  wire  T_7816;
  wire  T_7817;
  wire [63:0] T_7818;
  wire [63:0] GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire [1:0] GEN_127;
  wire [1:0] GEN_128;
  wire [2:0] GEN_129;
  wire  GEN_130;
  wire [3:0] GEN_131;
  wire  GEN_132;
  wire [4:0] GEN_133;
  wire [2:0] GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire [2:0] GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire [63:0] GEN_145;
  wire [63:0] GEN_146;
  wire [31:0] GEN_147;
  wire [39:0] GEN_148;
  wire  T_7819;
  wire  wb_set_sboard;
  wire  replay_wb_common;
  wire  T_7822;
  wire  T_7823;
  wire  replay_wb;
  wire  wb_xcpt;
  wire  T_7824;
  wire  T_7825;
  wire  T_7826;
  wire  dmem_resp_xpu;
  wire [7:0] dmem_resp_waddr;
  wire  dmem_resp_valid;
  wire  dmem_resp_replay;
  wire  T_7830;
  wire  T_7832;
  wire [63:0] ll_wdata;
  wire [7:0] ll_waddr;
  wire  T_7833;
  wire  ll_wen;
  wire  T_7834;
  wire  GEN_149;
  wire [7:0] GEN_150;
  wire  GEN_151;
  wire  T_7838;
  wire  T_7839;
  wire  T_7841;
  wire  wb_valid;
  wire  wb_wen;
  wire  rf_wen;
  wire [7:0] rf_waddr;
  wire  T_7842;
  wire  T_7843;
  wire [63:0] T_7844;
  wire [63:0] T_7845;
  wire [63:0] rf_wdata;
  wire [7:0] GEN_195;
  wire  T_7847;
  wire [4:0] T_7848;
  wire [4:0] T_7849;
  wire [7:0] GEN_196;
  wire  T_7851;
  wire [63:0] GEN_152;
  wire [7:0] GEN_197;
  wire  T_7852;
  wire [63:0] GEN_153;
  wire [63:0] GEN_159;
  wire [63:0] GEN_160;
  wire  GEN_163;
  wire [63:0] GEN_166;
  wire [63:0] GEN_167;
  wire [25:0] T_7853;
  wire [1:0] T_7854;
  wire [1:0] T_7855;
  wire  T_7857;
  wire  T_7859;
  wire  T_7860;
  wire  T_7862;
  wire [25:0] T_7863;
  wire  T_7865;
  wire  T_7868;
  wire  T_7869;
  wire  T_7871;
  wire  T_7872;
  wire  T_7873;
  wire  T_7874;
  wire [38:0] T_7875;
  wire [39:0] T_7876;
  wire [39:0] T_7877;
  wire [11:0] T_7894;
  wire [2:0] T_7895;
  wire  T_7897;
  wire  T_7898;
  wire  T_7900;
  wire  T_7901;
  wire  T_7903;
  wire  T_7904;
  reg [31:0] T_7906;
  reg [31:0] GEN_423;
  wire [255:0] GEN_211;
  wire [255:0] T_7909;
  wire [255:0] T_7911;
  wire [255:0] T_7912;
  wire [255:0] GEN_212;
  wire [255:0] T_7913;
  wire [255:0] GEN_168;
  wire [31:0] T_7915;
  wire  T_7916;
  wire  T_7917;
  wire [31:0] T_7918;
  wire  T_7919;
  wire  T_7920;
  wire [31:0] T_7921;
  wire  T_7922;
  wire  T_7923;
  wire  T_7924;
  wire  id_sboard_hazard;
  wire  T_7925;
  wire [31:0] GEN_213;
  wire [31:0] T_7927;
  wire [31:0] T_7929;
  wire [255:0] GEN_214;
  wire [255:0] T_7930;
  wire  T_7931;
  wire [255:0] GEN_169;
  wire  T_7932;
  wire  T_7933;
  wire  T_7934;
  wire  T_7935;
  wire  T_7936;
  wire  ex_cannot_bypass;
  wire  T_7937;
  wire  T_7938;
  wire  T_7939;
  wire  T_7940;
  wire  T_7941;
  wire  T_7942;
  wire  T_7943;
  wire  T_7944;
  wire  data_hazard_ex;
  wire  T_7946;
  wire  T_7948;
  wire  T_7949;
  wire  T_7950;
  wire  T_7952;
  wire  T_7953;
  wire  T_7954;
  wire  T_7955;
  wire  fp_data_hazard_ex;
  wire  T_7956;
  wire  T_7957;
  wire  id_ex_hazard;
  wire  T_7959;
  wire  T_7960;
  wire  T_7961;
  wire  T_7962;
  wire  T_7963;
  wire  mem_cannot_bypass;
  wire  T_7964;
  wire  T_7965;
  wire  T_7966;
  wire  T_7967;
  wire  T_7968;
  wire  T_7969;
  wire  T_7970;
  wire  T_7971;
  wire  data_hazard_mem;
  wire  T_7973;
  wire  T_7975;
  wire  T_7976;
  wire  T_7977;
  wire  T_7979;
  wire  T_7980;
  wire  T_7981;
  wire  T_7982;
  wire  fp_data_hazard_mem;
  wire  T_7983;
  wire  T_7984;
  wire  id_mem_hazard;
  wire  T_7985;
  wire  T_7986;
  wire  T_7987;
  wire  T_7988;
  wire  T_7989;
  wire  T_7990;
  wire  T_7991;
  wire  T_7992;
  wire  T_7993;
  wire  T_7994;
  wire  data_hazard_wb;
  wire  T_7996;
  wire  T_7998;
  wire  T_7999;
  wire  T_8000;
  wire  T_8002;
  wire  T_8003;
  wire  T_8004;
  wire  T_8005;
  wire  fp_data_hazard_wb;
  wire  T_8006;
  wire  T_8007;
  wire  id_wb_hazard;
  reg  dcache_blocked;
  reg [31:0] GEN_424;
  wire  T_8011;
  wire  T_8012;
  reg  rocc_blocked;
  reg [31:0] GEN_425;
  wire  T_8015;
  wire  T_8018;
  wire  T_8019;
  wire  T_8020;
  wire  T_8021;
  wire  T_8022;
  wire  T_8023;
  wire  T_8026;
  wire  T_8027;
  wire  T_8028;
  wire  T_8029;
  wire  T_8030;
  wire  ctrl_stalld;
  wire  T_8032;
  wire  T_8033;
  wire  T_8034;
  wire  T_8035;
  wire  T_8036;
  wire [39:0] T_8037;
  wire [39:0] T_8038;
  wire  T_8039;
  wire  T_8041;
  wire  T_8042;
  wire  T_8044;
  wire  T_8045;
  wire  T_8046;
  wire  T_8049;
  wire  T_8050;
  wire  T_8051;
  wire  T_8054;
  wire  T_8055;
  wire [4:0] T_8056;
  wire [4:0] T_8059;
  wire [4:0] GEN_215;
  wire  T_8060;
  wire  T_8061;
  wire  T_8062;
  wire  T_8065;
  wire  T_8066;
  wire  T_8069;
  wire  T_8072;
  wire  T_8073;
  wire  T_8074;
  wire  T_8077;
  wire  T_8078;
  wire  T_8079;
  wire [5:0] ex_dcache_tag;
  wire [25:0] T_8081;
  wire [1:0] T_8082;
  wire [1:0] T_8083;
  wire  T_8085;
  wire  T_8087;
  wire  T_8088;
  wire  T_8090;
  wire [25:0] T_8091;
  wire  T_8093;
  wire  T_8096;
  wire  T_8097;
  wire  T_8099;
  wire  T_8100;
  wire  T_8101;
  wire  T_8102;
  wire [38:0] T_8103;
  wire [39:0] T_8104;
  wire [63:0] T_8106;
  wire  T_8109;
  wire  T_8110;
  wire  T_8113;
  wire [6:0] T_8132_funct;
  wire [4:0] T_8132_rs2;
  wire [4:0] T_8132_rs1;
  wire  T_8132_xd;
  wire  T_8132_xs1;
  wire  T_8132_xs2;
  wire [4:0] T_8132_rd;
  wire [6:0] T_8132_opcode;
  wire [31:0] T_8142;
  wire [6:0] T_8143;
  wire [4:0] T_8144;
  wire  T_8145;
  wire  T_8146;
  wire  T_8147;
  wire [4:0] T_8148;
  wire [4:0] T_8149;
  wire [6:0] T_8150;
  wire [31:0] T_8151;
  wire [7:0] T_8153;
  wire [4:0] T_8154;
  reg [63:0] T_8155;
  reg [63:0] GEN_426;
  reg [63:0] T_8156;
  reg [63:0] GEN_427;
  wire [4:0] T_8157;
  reg [63:0] T_8158;
  reg [63:0] GEN_428;
  reg [63:0] T_8159;
  reg [63:0] GEN_429;
  wire  T_8161;
  reg  GEN_154;
  reg [31:0] GEN_430;
  reg [63:0] GEN_155;
  reg [63:0] GEN_431;
  reg  GEN_156;
  reg [31:0] GEN_432;
  reg [4:0] GEN_157;
  reg [31:0] GEN_433;
  reg  GEN_158;
  reg [31:0] GEN_434;
  reg  GEN_161;
  reg [31:0] GEN_435;
  reg  GEN_162;
  reg [31:0] GEN_436;
  reg  GEN_164;
  reg [31:0] GEN_437;
  reg  GEN_165;
  reg [31:0] GEN_438;
  reg  GEN_171;
  reg [31:0] GEN_439;
  reg  GEN_172;
  reg [31:0] GEN_440;
  reg  GEN_174;
  reg [31:0] GEN_441;
  reg  GEN_175;
  reg [31:0] GEN_442;
  reg  GEN_176;
  reg [31:0] GEN_443;
  reg  GEN_178;
  reg [31:0] GEN_444;
  reg  GEN_180;
  reg [31:0] GEN_445;
  reg  GEN_185;
  reg [31:0] GEN_446;
  reg  GEN_191;
  reg [31:0] GEN_447;
  reg  GEN_193;
  reg [31:0] GEN_448;
  reg  GEN_198;
  reg [31:0] GEN_449;
  reg [2:0] GEN_199;
  reg [31:0] GEN_450;
  reg [1:0] GEN_200;
  reg [31:0] GEN_451;
  reg [64:0] GEN_201;
  reg [95:0] GEN_452;
  reg [64:0] GEN_202;
  reg [95:0] GEN_453;
  reg [64:0] GEN_203;
  reg [95:0] GEN_454;
  reg  GEN_204;
  reg [31:0] GEN_455;
  reg  GEN_205;
  reg [31:0] GEN_456;
  reg  GEN_206;
  reg [31:0] GEN_457;
  reg  GEN_207;
  reg [31:0] GEN_458;
  reg  GEN_208;
  reg [31:0] GEN_459;
  reg [39:0] GEN_209;
  reg [63:0] GEN_460;
  reg [8:0] GEN_210;
  reg [31:0] GEN_461;
  reg [4:0] GEN_216;
  reg [31:0] GEN_462;
  reg [2:0] GEN_217;
  reg [31:0] GEN_463;
  reg [63:0] GEN_218;
  reg [63:0] GEN_464;
  reg  GEN_219;
  reg [31:0] GEN_465;
  reg  GEN_220;
  reg [31:0] GEN_466;
  reg [63:0] GEN_221;
  reg [63:0] GEN_467;
  reg [63:0] GEN_222;
  reg [63:0] GEN_468;
  reg  GEN_223;
  reg [31:0] GEN_469;
  reg  GEN_224;
  reg [31:0] GEN_470;
  reg  GEN_225;
  reg [31:0] GEN_471;
  reg  GEN_226;
  reg [31:0] GEN_472;
  reg  GEN_227;
  reg [31:0] GEN_473;
  reg  GEN_228;
  reg [31:0] GEN_474;
  reg  GEN_229;
  reg [31:0] GEN_475;
  reg  GEN_230;
  reg [31:0] GEN_476;
  reg [2:0] GEN_231;
  reg [31:0] GEN_477;
  reg [1:0] GEN_232;
  reg [31:0] GEN_478;
  reg [2:0] GEN_233;
  reg [31:0] GEN_479;
  reg  GEN_234;
  reg [31:0] GEN_480;
  reg [3:0] GEN_235;
  reg [31:0] GEN_481;
  reg [63:0] GEN_236;
  reg [63:0] GEN_482;
  reg  GEN_237;
  reg [31:0] GEN_483;
  reg  GEN_238;
  reg [31:0] GEN_484;
  reg [64:0] GEN_239;
  reg [95:0] GEN_485;
  reg [4:0] GEN_240;
  reg [31:0] GEN_486;
  reg  GEN_241;
  reg [31:0] GEN_487;
  reg  GEN_242;
  reg [31:0] GEN_488;
  reg  GEN_243;
  reg [31:0] GEN_489;
  reg [4:0] GEN_244;
  reg [31:0] GEN_490;
  reg [63:0] GEN_245;
  reg [63:0] GEN_491;
  reg  GEN_246;
  reg [31:0] GEN_492;
  reg [39:0] GEN_247;
  reg [63:0] GEN_493;
  reg [8:0] GEN_248;
  reg [31:0] GEN_494;
  reg [4:0] GEN_249;
  reg [31:0] GEN_495;
  reg [2:0] GEN_250;
  reg [31:0] GEN_496;
  reg  GEN_251;
  reg [31:0] GEN_497;
  reg [63:0] GEN_252;
  reg [63:0] GEN_498;
  reg  GEN_253;
  reg [31:0] GEN_499;
  reg [63:0] GEN_254;
  reg [63:0] GEN_500;
  reg  GEN_255;
  reg [31:0] GEN_501;
  reg  GEN_256;
  reg [31:0] GEN_502;
  reg  GEN_257;
  reg [31:0] GEN_503;
  reg [25:0] GEN_258;
  reg [31:0] GEN_504;
  reg [1:0] GEN_259;
  reg [31:0] GEN_505;
  reg [2:0] GEN_260;
  reg [31:0] GEN_506;
  reg  GEN_261;
  reg [31:0] GEN_507;
  reg [2:0] GEN_262;
  reg [31:0] GEN_508;
  reg [11:0] GEN_263;
  reg [31:0] GEN_509;
  reg [63:0] GEN_264;
  reg [63:0] GEN_510;
  reg  GEN_265;
  reg [31:0] GEN_511;
  reg  GEN_266;
  reg [31:0] GEN_512;
  reg [4:0] GEN_267;
  reg [31:0] GEN_513;
  reg  GEN_268;
  reg [31:0] GEN_514;
  reg  GEN_269;
  reg [31:0] GEN_515;
  reg  GEN_270;
  reg [31:0] GEN_516;
  reg  GEN_271;
  reg [31:0] GEN_517;
  reg  GEN_272;
  reg [31:0] GEN_518;
  reg  GEN_273;
  reg [31:0] GEN_519;
  reg  GEN_274;
  reg [31:0] GEN_520;
  reg  GEN_275;
  reg [31:0] GEN_521;
  reg  GEN_276;
  reg [31:0] GEN_522;
  reg  GEN_277;
  reg [31:0] GEN_523;
  reg  GEN_278;
  reg [31:0] GEN_524;
  reg  GEN_279;
  reg [31:0] GEN_525;
  reg  GEN_280;
  reg [31:0] GEN_526;
  reg  GEN_281;
  reg [31:0] GEN_527;
  reg  GEN_282;
  reg [31:0] GEN_528;
  reg  GEN_283;
  reg [31:0] GEN_529;
  reg [2:0] GEN_284;
  reg [31:0] GEN_530;
  reg [1:0] GEN_285;
  reg [31:0] GEN_531;
  reg [64:0] GEN_286;
  reg [95:0] GEN_532;
  reg [64:0] GEN_287;
  reg [95:0] GEN_533;
  reg [64:0] GEN_288;
  reg [95:0] GEN_534;
  reg  GEN_289;
  reg [31:0] GEN_535;
  CSRFile csr (
    .clk(csr_clk),
    .reset(csr_reset),
    .io_prci_reset(csr_io_prci_reset),
    .io_prci_id(csr_io_prci_id),
    .io_prci_interrupts_meip(csr_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(csr_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(csr_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(csr_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(csr_io_prci_interrupts_msip),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_csr_stall(csr_io_csr_stall),
    .io_csr_xcpt(csr_io_csr_xcpt),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero3(csr_io_status_zero3),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_vm(csr_io_status_vm),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_pum(csr_io_status_pum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_asid(csr_io_ptbr_asid),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_uarch_counters_0(csr_io_uarch_counters_0),
    .io_uarch_counters_1(csr_io_uarch_counters_1),
    .io_uarch_counters_2(csr_io_uarch_counters_2),
    .io_uarch_counters_3(csr_io_uarch_counters_3),
    .io_uarch_counters_4(csr_io_uarch_counters_4),
    .io_uarch_counters_5(csr_io_uarch_counters_5),
    .io_uarch_counters_6(csr_io_uarch_counters_6),
    .io_uarch_counters_7(csr_io_uarch_counters_7),
    .io_uarch_counters_8(csr_io_uarch_counters_8),
    .io_uarch_counters_9(csr_io_uarch_counters_9),
    .io_uarch_counters_10(csr_io_uarch_counters_10),
    .io_uarch_counters_11(csr_io_uarch_counters_11),
    .io_uarch_counters_12(csr_io_uarch_counters_12),
    .io_uarch_counters_13(csr_io_uarch_counters_13),
    .io_uarch_counters_14(csr_io_uarch_counters_14),
    .io_uarch_counters_15(csr_io_uarch_counters_15),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_badaddr(csr_io_badaddr),
    .io_fatc(csr_io_fatc),
    .io_time(csr_io_time),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_rocc_cmd_ready(csr_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(csr_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(csr_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(csr_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(csr_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(csr_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(csr_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(csr_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(csr_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(csr_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(csr_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(csr_io_rocc_cmd_bits_rs2),
    .io_rocc_resp_ready(csr_io_rocc_resp_ready),
    .io_rocc_resp_valid(csr_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(csr_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(csr_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(csr_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(csr_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(csr_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(csr_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(csr_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(csr_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(csr_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(csr_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(csr_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(csr_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(csr_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(csr_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(csr_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(csr_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(csr_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(csr_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(csr_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(csr_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(csr_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(csr_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(csr_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(csr_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(csr_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(csr_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(csr_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(csr_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(csr_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(csr_io_rocc_mem_ordered),
    .io_rocc_busy(csr_io_rocc_busy),
    .io_rocc_status_debug(csr_io_rocc_status_debug),
    .io_rocc_status_prv(csr_io_rocc_status_prv),
    .io_rocc_status_sd(csr_io_rocc_status_sd),
    .io_rocc_status_zero3(csr_io_rocc_status_zero3),
    .io_rocc_status_sd_rv32(csr_io_rocc_status_sd_rv32),
    .io_rocc_status_zero2(csr_io_rocc_status_zero2),
    .io_rocc_status_vm(csr_io_rocc_status_vm),
    .io_rocc_status_zero1(csr_io_rocc_status_zero1),
    .io_rocc_status_pum(csr_io_rocc_status_pum),
    .io_rocc_status_mprv(csr_io_rocc_status_mprv),
    .io_rocc_status_xs(csr_io_rocc_status_xs),
    .io_rocc_status_fs(csr_io_rocc_status_fs),
    .io_rocc_status_mpp(csr_io_rocc_status_mpp),
    .io_rocc_status_hpp(csr_io_rocc_status_hpp),
    .io_rocc_status_spp(csr_io_rocc_status_spp),
    .io_rocc_status_mpie(csr_io_rocc_status_mpie),
    .io_rocc_status_hpie(csr_io_rocc_status_hpie),
    .io_rocc_status_spie(csr_io_rocc_status_spie),
    .io_rocc_status_upie(csr_io_rocc_status_upie),
    .io_rocc_status_mie(csr_io_rocc_status_mie),
    .io_rocc_status_hie(csr_io_rocc_status_hie),
    .io_rocc_status_sie(csr_io_rocc_status_sie),
    .io_rocc_status_uie(csr_io_rocc_status_uie),
    .io_rocc_interrupt(csr_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(csr_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(csr_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(csr_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(csr_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(csr_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(csr_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(csr_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(csr_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(csr_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(csr_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(csr_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(csr_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(csr_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(csr_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(csr_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(csr_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(csr_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(csr_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(csr_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(csr_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(csr_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(csr_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(csr_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(csr_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(csr_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(csr_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(csr_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(csr_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(csr_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(csr_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(csr_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(csr_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(csr_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(csr_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(csr_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(csr_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(csr_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(csr_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(csr_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(csr_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(csr_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(csr_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(csr_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(csr_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(csr_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(csr_io_rocc_exception),
    .io_rocc_csr_waddr(csr_io_rocc_csr_waddr),
    .io_rocc_csr_wdata(csr_io_rocc_csr_wdata),
    .io_rocc_csr_wen(csr_io_rocc_csr_wen),
    .io_rocc_host_id(csr_io_rocc_host_id),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_tdrtype(csr_io_bp_0_control_tdrtype),
    .io_bp_0_control_bpamaskmax(csr_io_bp_0_control_bpamaskmax),
    .io_bp_0_control_reserved(csr_io_bp_0_control_reserved),
    .io_bp_0_control_bpaction(csr_io_bp_0_control_bpaction),
    .io_bp_0_control_bpmatch(csr_io_bp_0_control_bpmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_h(csr_io_bp_0_control_h),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_address(csr_io_bp_0_address)
  );
  BreakpointUnit bpu (
    .clk(bpu_clk),
    .reset(bpu_reset),
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_status_sd(bpu_io_status_sd),
    .io_status_zero3(bpu_io_status_zero3),
    .io_status_sd_rv32(bpu_io_status_sd_rv32),
    .io_status_zero2(bpu_io_status_zero2),
    .io_status_vm(bpu_io_status_vm),
    .io_status_zero1(bpu_io_status_zero1),
    .io_status_pum(bpu_io_status_pum),
    .io_status_mprv(bpu_io_status_mprv),
    .io_status_xs(bpu_io_status_xs),
    .io_status_fs(bpu_io_status_fs),
    .io_status_mpp(bpu_io_status_mpp),
    .io_status_hpp(bpu_io_status_hpp),
    .io_status_spp(bpu_io_status_spp),
    .io_status_mpie(bpu_io_status_mpie),
    .io_status_hpie(bpu_io_status_hpie),
    .io_status_spie(bpu_io_status_spie),
    .io_status_upie(bpu_io_status_upie),
    .io_status_mie(bpu_io_status_mie),
    .io_status_hie(bpu_io_status_hie),
    .io_status_sie(bpu_io_status_sie),
    .io_status_uie(bpu_io_status_uie),
    .io_bp_0_control_tdrtype(bpu_io_bp_0_control_tdrtype),
    .io_bp_0_control_bpamaskmax(bpu_io_bp_0_control_bpamaskmax),
    .io_bp_0_control_reserved(bpu_io_bp_0_control_reserved),
    .io_bp_0_control_bpaction(bpu_io_bp_0_control_bpaction),
    .io_bp_0_control_bpmatch(bpu_io_bp_0_control_bpmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_h(bpu_io_bp_0_control_h),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st)
  );
  ALU alu (
    .clk(alu_clk),
    .reset(alu_reset),
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  MulDiv div (
    .clk(div_clk),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag)
  );
  assign io_imem_req_valid = take_pc_mem_wb;
  assign io_imem_req_bits_pc = T_8038;
  assign io_imem_resp_ready = T_8046;
  assign io_imem_btb_update_valid = T_8054;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign io_imem_btb_update_bits_pc = mem_reg_pc[38:0];
  assign io_imem_btb_update_bits_target = io_imem_req_bits_pc[38:0];
  assign io_imem_btb_update_bits_taken = GEN_154;
  assign io_imem_btb_update_bits_isJump = T_8055;
  assign io_imem_btb_update_bits_isReturn = T_8061;
  assign io_imem_btb_update_bits_br_pc = mem_reg_pc[38:0];
  assign io_imem_bht_update_valid = T_8065;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_pc = mem_reg_pc[38:0];
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_ras_update_valid = T_8072;
  assign io_imem_ras_update_bits_isCall = T_8074;
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_returnAddr = mem_int_wdata[38:0];
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_flush_icache = T_8042;
  assign io_imem_flush_tlb = csr_io_fatc;
  assign io_dmem_req_valid = T_8079;
  assign io_dmem_req_bits_addr = T_8104;
  assign io_dmem_req_bits_tag = {{3'd0}, ex_dcache_tag};
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_data = GEN_155;
  assign io_dmem_s1_kill = T_7801;
  assign io_dmem_s1_data = T_8106;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_ptw_ptbr_asid = csr_io_ptbr_asid;
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn;
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_status_debug = csr_io_status_debug;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_status_zero3 = csr_io_status_zero3;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_pum = csr_io_status_pum;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_mpp = csr_io_status_mpp;
  assign io_ptw_status_hpp = csr_io_status_hpp;
  assign io_ptw_status_spp = csr_io_status_spp;
  assign io_ptw_status_mpie = csr_io_status_mpie;
  assign io_ptw_status_hpie = csr_io_status_hpie;
  assign io_ptw_status_spie = csr_io_status_spie;
  assign io_ptw_status_upie = csr_io_status_upie;
  assign io_ptw_status_mie = csr_io_status_mie;
  assign io_ptw_status_hie = csr_io_status_hie;
  assign io_ptw_status_sie = csr_io_status_sie;
  assign io_ptw_status_uie = csr_io_status_uie;
  assign io_fpu_inst = io_imem_resp_bits_data_0;
  assign io_fpu_fromint_data = T_7375;
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_dmem_resp_val = T_8078;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr[4:0];
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
  assign io_fpu_valid = T_8077;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_killm = killm_common;
  assign io_fpu_cp_req_valid = GEN_156;
  assign io_fpu_cp_req_bits_cmd = GEN_157;
  assign io_fpu_cp_req_bits_ldst = GEN_158;
  assign io_fpu_cp_req_bits_wen = GEN_161;
  assign io_fpu_cp_req_bits_ren1 = GEN_162;
  assign io_fpu_cp_req_bits_ren2 = GEN_164;
  assign io_fpu_cp_req_bits_ren3 = GEN_165;
  assign io_fpu_cp_req_bits_swap12 = GEN_171;
  assign io_fpu_cp_req_bits_swap23 = GEN_172;
  assign io_fpu_cp_req_bits_single = GEN_174;
  assign io_fpu_cp_req_bits_fromint = GEN_175;
  assign io_fpu_cp_req_bits_toint = GEN_176;
  assign io_fpu_cp_req_bits_fastpipe = GEN_178;
  assign io_fpu_cp_req_bits_fma = GEN_180;
  assign io_fpu_cp_req_bits_div = GEN_185;
  assign io_fpu_cp_req_bits_sqrt = GEN_191;
  assign io_fpu_cp_req_bits_round = GEN_193;
  assign io_fpu_cp_req_bits_wflags = GEN_198;
  assign io_fpu_cp_req_bits_rm = GEN_199;
  assign io_fpu_cp_req_bits_typ = GEN_200;
  assign io_fpu_cp_req_bits_in1 = GEN_201;
  assign io_fpu_cp_req_bits_in2 = GEN_202;
  assign io_fpu_cp_req_bits_in3 = GEN_203;
  assign io_fpu_cp_resp_ready = GEN_204;
  assign io_rocc_cmd_valid = T_8110;
  assign io_rocc_cmd_bits_inst_funct = T_8132_funct;
  assign io_rocc_cmd_bits_inst_rs2 = T_8132_rs2;
  assign io_rocc_cmd_bits_inst_rs1 = T_8132_rs1;
  assign io_rocc_cmd_bits_inst_xd = T_8132_xd;
  assign io_rocc_cmd_bits_inst_xs1 = T_8132_xs1;
  assign io_rocc_cmd_bits_inst_xs2 = T_8132_xs2;
  assign io_rocc_cmd_bits_inst_rd = T_8132_rd;
  assign io_rocc_cmd_bits_inst_opcode = T_8132_opcode;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign io_rocc_resp_ready = GEN_205;
  assign io_rocc_mem_req_ready = GEN_206;
  assign io_rocc_mem_s2_nack = GEN_207;
  assign io_rocc_mem_resp_valid = GEN_208;
  assign io_rocc_mem_resp_bits_addr = GEN_209;
  assign io_rocc_mem_resp_bits_tag = GEN_210;
  assign io_rocc_mem_resp_bits_cmd = GEN_216;
  assign io_rocc_mem_resp_bits_typ = GEN_217;
  assign io_rocc_mem_resp_bits_data = GEN_218;
  assign io_rocc_mem_resp_bits_replay = GEN_219;
  assign io_rocc_mem_resp_bits_has_data = GEN_220;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_221;
  assign io_rocc_mem_resp_bits_store_data = GEN_222;
  assign io_rocc_mem_replay_next = GEN_223;
  assign io_rocc_mem_xcpt_ma_ld = GEN_224;
  assign io_rocc_mem_xcpt_ma_st = GEN_225;
  assign io_rocc_mem_xcpt_pf_ld = GEN_226;
  assign io_rocc_mem_xcpt_pf_st = GEN_227;
  assign io_rocc_mem_ordered = GEN_228;
  assign io_rocc_status_debug = csr_io_status_debug;
  assign io_rocc_status_prv = csr_io_status_prv;
  assign io_rocc_status_sd = csr_io_status_sd;
  assign io_rocc_status_zero3 = csr_io_status_zero3;
  assign io_rocc_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_rocc_status_zero2 = csr_io_status_zero2;
  assign io_rocc_status_vm = csr_io_status_vm;
  assign io_rocc_status_zero1 = csr_io_status_zero1;
  assign io_rocc_status_pum = csr_io_status_pum;
  assign io_rocc_status_mprv = csr_io_status_mprv;
  assign io_rocc_status_xs = csr_io_status_xs;
  assign io_rocc_status_fs = csr_io_status_fs;
  assign io_rocc_status_mpp = csr_io_status_mpp;
  assign io_rocc_status_hpp = csr_io_status_hpp;
  assign io_rocc_status_spp = csr_io_status_spp;
  assign io_rocc_status_mpie = csr_io_status_mpie;
  assign io_rocc_status_hpie = csr_io_status_hpie;
  assign io_rocc_status_spie = csr_io_status_spie;
  assign io_rocc_status_upie = csr_io_status_upie;
  assign io_rocc_status_mie = csr_io_status_mie;
  assign io_rocc_status_hie = csr_io_status_hie;
  assign io_rocc_status_sie = csr_io_status_sie;
  assign io_rocc_status_uie = csr_io_status_uie;
  assign io_rocc_autl_acquire_ready = GEN_229;
  assign io_rocc_autl_grant_valid = GEN_230;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_231;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_232;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_233;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_234;
  assign io_rocc_autl_grant_bits_g_type = GEN_235;
  assign io_rocc_autl_grant_bits_data = GEN_236;
  assign io_rocc_fpu_req_ready = GEN_237;
  assign io_rocc_fpu_resp_valid = GEN_238;
  assign io_rocc_fpu_resp_bits_data = GEN_239;
  assign io_rocc_fpu_resp_bits_exc = GEN_240;
  assign io_rocc_exception = T_8113;
  assign io_rocc_csr_waddr = csr_io_rocc_csr_waddr;
  assign io_rocc_csr_wdata = csr_io_rocc_csr_wdata;
  assign io_rocc_csr_wen = csr_io_rocc_csr_wen;
  assign io_rocc_host_id = GEN_241;
  assign take_pc_mem = T_7733;
  assign take_pc_wb = T_7825;
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem;
  assign id_ctrl_legal = T_6769;
  assign id_ctrl_fp = 1'h0;
  assign id_ctrl_rocc = 1'h0;
  assign id_ctrl_branch = T_6775;
  assign id_ctrl_jal = T_6781;
  assign id_ctrl_jalr = T_6787;
  assign id_ctrl_rxs2 = T_6805;
  assign id_ctrl_rxs1 = T_6826;
  assign id_ctrl_sel_alu2 = T_6862;
  assign id_ctrl_sel_alu1 = T_6879;
  assign id_ctrl_sel_imm = T_6911;
  assign id_ctrl_alu_dw = T_6922;
  assign id_ctrl_alu_fn = T_7006;
  assign id_ctrl_mem = T_7022;
  assign id_ctrl_mem_cmd = T_7082;
  assign id_ctrl_mem_type = T_7102;
  assign id_ctrl_rfs1 = 1'h0;
  assign id_ctrl_rfs2 = 1'h0;
  assign id_ctrl_rfs3 = 1'h0;
  assign id_ctrl_wfd = 1'h0;
  assign id_ctrl_div = T_7110;
  assign id_ctrl_wxd = T_7140;
  assign id_ctrl_csr = T_7160;
  assign id_ctrl_fence_i = T_7164;
  assign id_ctrl_fence = T_7170;
  assign id_ctrl_amo = T_7176;
  assign T_6629 = io_imem_resp_bits_data_0 & 32'h405f;
  assign T_6631 = T_6629 == 32'h3;
  assign T_6633 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T_6635 = T_6633 == 32'h3;
  assign T_6637 = io_imem_resp_bits_data_0 & 32'h106f;
  assign T_6639 = T_6637 == 32'h3;
  assign T_6641 = io_imem_resp_bits_data_0 & 32'h607f;
  assign T_6643 = T_6641 == 32'hf;
  assign T_6645 = io_imem_resp_bits_data_0 & 32'h7077;
  assign T_6647 = T_6645 == 32'h13;
  assign T_6649 = io_imem_resp_bits_data_0 & 32'h5f;
  assign T_6651 = T_6649 == 32'h17;
  assign T_6653 = io_imem_resp_bits_data_0 & 32'hfc00007f;
  assign T_6655 = T_6653 == 32'h33;
  assign T_6657 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T_6659 = T_6657 == 32'h33;
  assign T_6661 = io_imem_resp_bits_data_0 & 32'h707b;
  assign T_6663 = T_6661 == 32'h63;
  assign T_6665 = io_imem_resp_bits_data_0 & 32'h7f;
  assign T_6667 = T_6665 == 32'h6f;
  assign T_6669 = io_imem_resp_bits_data_0 & 32'hffefffff;
  assign T_6671 = T_6669 == 32'h73;
  assign T_6673 = io_imem_resp_bits_data_0 & 32'hfc00305f;
  assign T_6675 = T_6673 == 32'h1013;
  assign T_6677 = io_imem_resp_bits_data_0 & 32'hfe00305f;
  assign T_6679 = T_6677 == 32'h101b;
  assign T_6683 = T_6633 == 32'h2013;
  assign T_6685 = io_imem_resp_bits_data_0 & 32'h1800607f;
  assign T_6687 = T_6685 == 32'h202f;
  assign T_6691 = T_6633 == 32'h2073;
  assign T_6693 = io_imem_resp_bits_data_0 & 32'hbc00707f;
  assign T_6695 = T_6693 == 32'h5013;
  assign T_6697 = io_imem_resp_bits_data_0 & 32'hbe00705f;
  assign T_6699 = T_6697 == 32'h501b;
  assign T_6703 = T_6657 == 32'h5033;
  assign T_6705 = io_imem_resp_bits_data_0 & 32'hfe004077;
  assign T_6707 = T_6705 == 32'h2004033;
  assign T_6709 = io_imem_resp_bits_data_0 & 32'he800607f;
  assign T_6711 = T_6709 == 32'h800202f;
  assign T_6713 = io_imem_resp_bits_data_0 & 32'hf9f0607f;
  assign T_6715 = T_6713 == 32'h1000202f;
  assign T_6717 = io_imem_resp_bits_data_0 & 32'hdfffffff;
  assign T_6719 = T_6717 == 32'h10200073;
  assign T_6721 = io_imem_resp_bits_data_0 & 32'hfff07fff;
  assign T_6723 = T_6721 == 32'h10400073;
  assign T_6725 = io_imem_resp_bits_data_0 == 32'h10500073;
  assign T_6727 = io_imem_resp_bits_data_0 == 32'h7b200073;
  assign T_6729 = io_imem_resp_bits_data_0 & 32'h306f;
  assign T_6731 = T_6729 == 32'h1063;
  assign T_6733 = io_imem_resp_bits_data_0 & 32'h407f;
  assign T_6735 = T_6733 == 32'h4063;
  assign T_6737 = io_imem_resp_bits_data_0 & 32'hfc007077;
  assign T_6739 = T_6737 == 32'h33;
  assign T_6742 = T_6631 | T_6635;
  assign T_6743 = T_6742 | T_6639;
  assign T_6744 = T_6743 | T_6643;
  assign T_6745 = T_6744 | T_6647;
  assign T_6746 = T_6745 | T_6651;
  assign T_6747 = T_6746 | T_6655;
  assign T_6748 = T_6747 | T_6659;
  assign T_6749 = T_6748 | T_6663;
  assign T_6750 = T_6749 | T_6667;
  assign T_6751 = T_6750 | T_6671;
  assign T_6752 = T_6751 | T_6675;
  assign T_6753 = T_6752 | T_6679;
  assign T_6754 = T_6753 | T_6683;
  assign T_6755 = T_6754 | T_6687;
  assign T_6756 = T_6755 | T_6691;
  assign T_6757 = T_6756 | T_6695;
  assign T_6758 = T_6757 | T_6699;
  assign T_6759 = T_6758 | T_6703;
  assign T_6760 = T_6759 | T_6707;
  assign T_6761 = T_6760 | T_6711;
  assign T_6762 = T_6761 | T_6715;
  assign T_6763 = T_6762 | T_6719;
  assign T_6764 = T_6763 | T_6723;
  assign T_6765 = T_6764 | T_6725;
  assign T_6766 = T_6765 | T_6727;
  assign T_6767 = T_6766 | T_6731;
  assign T_6768 = T_6767 | T_6735;
  assign T_6769 = T_6768 | T_6739;
  assign T_6773 = io_imem_resp_bits_data_0 & 32'h54;
  assign T_6775 = T_6773 == 32'h40;
  assign T_6779 = io_imem_resp_bits_data_0 & 32'h48;
  assign T_6781 = T_6779 == 32'h48;
  assign T_6785 = io_imem_resp_bits_data_0 & 32'h1c;
  assign T_6787 = T_6785 == 32'h4;
  assign T_6791 = io_imem_resp_bits_data_0 & 32'h70;
  assign T_6793 = T_6791 == 32'h20;
  assign T_6795 = io_imem_resp_bits_data_0 & 32'h64;
  assign T_6797 = T_6795 == 32'h20;
  assign T_6799 = io_imem_resp_bits_data_0 & 32'h34;
  assign T_6801 = T_6799 == 32'h20;
  assign T_6804 = T_6793 | T_6797;
  assign T_6805 = T_6804 | T_6801;
  assign T_6807 = io_imem_resp_bits_data_0 & 32'h4004;
  assign T_6809 = T_6807 == 32'h0;
  assign T_6811 = io_imem_resp_bits_data_0 & 32'h44;
  assign T_6813 = T_6811 == 32'h0;
  assign T_6815 = io_imem_resp_bits_data_0 & 32'h18;
  assign T_6817 = T_6815 == 32'h0;
  assign T_6819 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T_6821 = T_6819 == 32'h2000;
  assign T_6824 = T_6809 | T_6813;
  assign T_6825 = T_6824 | T_6817;
  assign T_6826 = T_6825 | T_6821;
  assign T_6828 = io_imem_resp_bits_data_0 & 32'h58;
  assign T_6830 = T_6828 == 32'h0;
  assign T_6832 = io_imem_resp_bits_data_0 & 32'h20;
  assign T_6834 = T_6832 == 32'h0;
  assign T_6836 = io_imem_resp_bits_data_0 & 32'hc;
  assign T_6838 = T_6836 == 32'h4;
  assign T_6840 = io_imem_resp_bits_data_0 & 32'h4050;
  assign T_6842 = T_6840 == 32'h4050;
  assign T_6845 = T_6830 | T_6834;
  assign T_6846 = T_6845 | T_6838;
  assign T_6847 = T_6846 | T_6781;
  assign T_6848 = T_6847 | T_6842;
  assign T_6852 = T_6779 == 32'h0;
  assign T_6854 = io_imem_resp_bits_data_0 & 32'h4008;
  assign T_6856 = T_6854 == 32'h4000;
  assign T_6859 = T_6852 | T_6813;
  assign T_6860 = T_6859 | T_6817;
  assign T_6861 = T_6860 | T_6856;
  assign T_6862 = {T_6861,T_6848};
  assign T_6864 = io_imem_resp_bits_data_0 & 32'h50;
  assign T_6866 = T_6864 == 32'h0;
  assign T_6869 = T_6809 | T_6866;
  assign T_6870 = T_6869 | T_6813;
  assign T_6871 = T_6870 | T_6817;
  assign T_6873 = io_imem_resp_bits_data_0 & 32'h24;
  assign T_6875 = T_6873 == 32'h4;
  assign T_6878 = T_6875 | T_6781;
  assign T_6879 = {T_6878,T_6871};
  assign T_6883 = T_6815 == 32'h8;
  assign T_6887 = T_6811 == 32'h40;
  assign T_6890 = T_6883 | T_6887;
  assign T_6894 = T_6811 == 32'h4;
  assign T_6897 = T_6894 | T_6883;
  assign T_6901 = T_6873 == 32'h0;
  assign T_6903 = io_imem_resp_bits_data_0 & 32'h14;
  assign T_6905 = T_6903 == 32'h10;
  assign T_6908 = T_6901 | T_6787;
  assign T_6909 = T_6908 | T_6905;
  assign T_6910 = {T_6897,T_6890};
  assign T_6911 = {T_6909,T_6910};
  assign T_6913 = io_imem_resp_bits_data_0 & 32'h10;
  assign T_6915 = T_6913 == 32'h0;
  assign T_6917 = io_imem_resp_bits_data_0 & 32'h8;
  assign T_6919 = T_6917 == 32'h0;
  assign T_6922 = T_6915 | T_6919;
  assign T_6924 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T_6926 = T_6924 == 32'h1010;
  assign T_6928 = io_imem_resp_bits_data_0 & 32'h1058;
  assign T_6930 = T_6928 == 32'h1040;
  assign T_6932 = io_imem_resp_bits_data_0 & 32'h7044;
  assign T_6934 = T_6932 == 32'h7000;
  assign T_6937 = T_6926 | T_6930;
  assign T_6938 = T_6937 | T_6934;
  assign T_6940 = io_imem_resp_bits_data_0 & 32'h4054;
  assign T_6942 = T_6940 == 32'h40;
  assign T_6944 = io_imem_resp_bits_data_0 & 32'h2058;
  assign T_6946 = T_6944 == 32'h2040;
  assign T_6950 = T_6924 == 32'h3010;
  assign T_6952 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T_6954 = T_6952 == 32'h6010;
  assign T_6956 = io_imem_resp_bits_data_0 & 32'h40003034;
  assign T_6958 = T_6956 == 32'h40000030;
  assign T_6960 = io_imem_resp_bits_data_0 & 32'h40001054;
  assign T_6962 = T_6960 == 32'h40001010;
  assign T_6965 = T_6942 | T_6946;
  assign T_6966 = T_6965 | T_6950;
  assign T_6967 = T_6966 | T_6954;
  assign T_6968 = T_6967 | T_6958;
  assign T_6969 = T_6968 | T_6962;
  assign T_6971 = io_imem_resp_bits_data_0 & 32'h2054;
  assign T_6973 = T_6971 == 32'h2010;
  assign T_6975 = io_imem_resp_bits_data_0 & 32'h40004054;
  assign T_6977 = T_6975 == 32'h4010;
  assign T_6979 = io_imem_resp_bits_data_0 & 32'h5054;
  assign T_6981 = T_6979 == 32'h4010;
  assign T_6983 = io_imem_resp_bits_data_0 & 32'h4058;
  assign T_6985 = T_6983 == 32'h4040;
  assign T_6988 = T_6973 | T_6977;
  assign T_6989 = T_6988 | T_6981;
  assign T_6990 = T_6989 | T_6985;
  assign T_6994 = T_6952 == 32'h2010;
  assign T_6996 = io_imem_resp_bits_data_0 & 32'h40003054;
  assign T_6998 = T_6996 == 32'h40001010;
  assign T_7001 = T_6994 | T_6985;
  assign T_7002 = T_7001 | T_6958;
  assign T_7003 = T_7002 | T_6998;
  assign T_7004 = {T_6969,T_6938};
  assign T_7005 = {T_6990,T_7004};
  assign T_7006 = {T_7003,T_7005};
  assign T_7008 = io_imem_resp_bits_data_0 & 32'h107f;
  assign T_7010 = T_7008 == 32'h3;
  assign T_7012 = io_imem_resp_bits_data_0 & 32'h707f;
  assign T_7014 = T_7012 == 32'h100f;
  assign T_7018 = T_6742 | T_7010;
  assign T_7019 = T_7018 | T_7014;
  assign T_7020 = T_7019 | T_6687;
  assign T_7021 = T_7020 | T_6711;
  assign T_7022 = T_7021 | T_6715;
  assign T_7024 = io_imem_resp_bits_data_0 & 32'h2008;
  assign T_7026 = T_7024 == 32'h8;
  assign T_7028 = io_imem_resp_bits_data_0 & 32'h28;
  assign T_7030 = T_7028 == 32'h20;
  assign T_7032 = io_imem_resp_bits_data_0 & 32'h18000020;
  assign T_7034 = T_7032 == 32'h18000020;
  assign T_7036 = io_imem_resp_bits_data_0 & 32'h20000020;
  assign T_7038 = T_7036 == 32'h20000020;
  assign T_7041 = T_7026 | T_7030;
  assign T_7042 = T_7041 | T_7034;
  assign T_7043 = T_7042 | T_7038;
  assign T_7045 = io_imem_resp_bits_data_0 & 32'h10002008;
  assign T_7047 = T_7045 == 32'h10002008;
  assign T_7049 = io_imem_resp_bits_data_0 & 32'h40002008;
  assign T_7051 = T_7049 == 32'h40002008;
  assign T_7054 = T_7047 | T_7051;
  assign T_7056 = io_imem_resp_bits_data_0 & 32'h8000008;
  assign T_7058 = T_7056 == 32'h8000008;
  assign T_7060 = io_imem_resp_bits_data_0 & 32'h10000008;
  assign T_7062 = T_7060 == 32'h10000008;
  assign T_7064 = io_imem_resp_bits_data_0 & 32'h80000008;
  assign T_7066 = T_7064 == 32'h80000008;
  assign T_7069 = T_7026 | T_7058;
  assign T_7070 = T_7069 | T_7062;
  assign T_7071 = T_7070 | T_7066;
  assign T_7073 = io_imem_resp_bits_data_0 & 32'h18002008;
  assign T_7075 = T_7073 == 32'h2008;
  assign T_7079 = {T_7054,T_7043};
  assign T_7080 = {T_7071,T_7079};
  assign T_7081 = {T_7075,T_7080};
  assign T_7082 = {1'h0,T_7081};
  assign T_7084 = io_imem_resp_bits_data_0 & 32'h1000;
  assign T_7086 = T_7084 == 32'h1000;
  assign T_7090 = io_imem_resp_bits_data_0 & 32'h2000;
  assign T_7092 = T_7090 == 32'h2000;
  assign T_7096 = io_imem_resp_bits_data_0 & 32'h4000;
  assign T_7098 = T_7096 == 32'h4000;
  assign T_7101 = {T_7092,T_7086};
  assign T_7102 = {T_7098,T_7101};
  assign T_7108 = io_imem_resp_bits_data_0 & 32'h2000074;
  assign T_7110 = T_7108 == 32'h2000030;
  assign T_7116 = T_6864 == 32'h10;
  assign T_7118 = io_imem_resp_bits_data_0 & 32'h1010;
  assign T_7120 = T_7118 == 32'h1010;
  assign T_7124 = T_7024 == 32'h2008;
  assign T_7126 = io_imem_resp_bits_data_0 & 32'h2010;
  assign T_7128 = T_7126 == 32'h2010;
  assign T_7132 = T_7028 == 32'h0;
  assign T_7135 = T_6838 | T_7116;
  assign T_7136 = T_7135 | T_6781;
  assign T_7137 = T_7136 | T_7120;
  assign T_7138 = T_7137 | T_7124;
  assign T_7139 = T_7138 | T_7128;
  assign T_7140 = T_7139 | T_7132;
  assign T_7142 = io_imem_resp_bits_data_0 & 32'h1050;
  assign T_7144 = T_7142 == 32'h1050;
  assign T_7150 = T_6819 == 32'h2050;
  assign T_7154 = io_imem_resp_bits_data_0 & 32'h3050;
  assign T_7156 = T_7154 == 32'h50;
  assign T_7159 = {T_7150,T_7144};
  assign T_7160 = {T_7156,T_7159};
  assign T_7162 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T_7164 = T_7162 == 32'h1008;
  assign T_7170 = T_7162 == 32'h8;
  assign T_7174 = io_imem_resp_bits_data_0 & 32'h6048;
  assign T_7176 = T_7174 == 32'h2008;
  assign id_raddr3 = io_imem_resp_bits_data_0[31:27];
  assign id_raddr2 = io_imem_resp_bits_data_0[24:20];
  assign id_raddr1 = io_imem_resp_bits_data_0[19:15];
  assign id_waddr = io_imem_resp_bits_data_0[11:7];
  assign id_load_use = T_7986;
  assign T_7183_T_7193_addr = T_7192;
  assign T_7183_T_7193_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_7183_T_7193_data = T_7183[T_7183_T_7193_addr];
  `else
  assign T_7183_T_7193_data = T_7183_T_7193_addr >= 5'h1f ? $random : T_7183[T_7183_T_7193_addr];
  `endif
  assign T_7183_T_7204_addr = T_7203;
  assign T_7183_T_7204_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_7183_T_7204_data = T_7183[T_7183_T_7204_addr];
  `else
  assign T_7183_T_7204_data = T_7183_T_7204_addr >= 5'h1f ? $random : T_7183[T_7183_T_7204_addr];
  `endif
  assign T_7183_T_7850_data = rf_wdata;
  assign T_7183_T_7850_addr = T_7849;
  assign T_7183_T_7850_mask = GEN_163;
  assign T_7183_T_7850_en = GEN_163;
  assign T_7185 = GEN_166;
  assign GEN_170 = {{4'd0}, 1'h0};
  assign T_7188 = id_raddr1 == GEN_170;
  assign T_7192 = ~ id_raddr1;
  assign T_7194 = T_7183_T_7193_data;
  assign T_7196 = GEN_167;
  assign T_7203 = ~ id_raddr2;
  assign T_7205 = T_7183_T_7204_data;
  assign ctrl_killd = T_8035;
  assign csr_clk = clk;
  assign csr_reset = reset;
  assign csr_io_prci_reset = io_prci_reset;
  assign csr_io_prci_id = io_prci_id;
  assign csr_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign csr_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign csr_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign csr_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign csr_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign csr_io_rw_addr = T_7894;
  assign csr_io_rw_cmd = T_7895;
  assign csr_io_rw_wdata = wb_reg_wdata;
  assign csr_io_exception = wb_reg_xcpt;
  assign csr_io_retire = wb_valid;
  assign csr_io_uarch_counters_0 = 1'h0;
  assign csr_io_uarch_counters_1 = 1'h0;
  assign csr_io_uarch_counters_2 = 1'h0;
  assign csr_io_uarch_counters_3 = 1'h0;
  assign csr_io_uarch_counters_4 = 1'h0;
  assign csr_io_uarch_counters_5 = 1'h0;
  assign csr_io_uarch_counters_6 = 1'h0;
  assign csr_io_uarch_counters_7 = 1'h0;
  assign csr_io_uarch_counters_8 = 1'h0;
  assign csr_io_uarch_counters_9 = 1'h0;
  assign csr_io_uarch_counters_10 = 1'h0;
  assign csr_io_uarch_counters_11 = 1'h0;
  assign csr_io_uarch_counters_12 = 1'h0;
  assign csr_io_uarch_counters_13 = 1'h0;
  assign csr_io_uarch_counters_14 = 1'h0;
  assign csr_io_uarch_counters_15 = 1'h0;
  assign csr_io_cause = wb_reg_cause;
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_badaddr = T_7877;
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid;
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits;
  assign csr_io_rocc_cmd_ready = GEN_242;
  assign csr_io_rocc_resp_valid = GEN_243;
  assign csr_io_rocc_resp_bits_rd = GEN_244;
  assign csr_io_rocc_resp_bits_data = GEN_245;
  assign csr_io_rocc_mem_req_valid = GEN_246;
  assign csr_io_rocc_mem_req_bits_addr = GEN_247;
  assign csr_io_rocc_mem_req_bits_tag = GEN_248;
  assign csr_io_rocc_mem_req_bits_cmd = GEN_249;
  assign csr_io_rocc_mem_req_bits_typ = GEN_250;
  assign csr_io_rocc_mem_req_bits_phys = GEN_251;
  assign csr_io_rocc_mem_req_bits_data = GEN_252;
  assign csr_io_rocc_mem_s1_kill = GEN_253;
  assign csr_io_rocc_mem_s1_data = GEN_254;
  assign csr_io_rocc_mem_invalidate_lr = GEN_255;
  assign csr_io_rocc_busy = GEN_256;
  assign csr_io_rocc_interrupt = io_rocc_interrupt;
  assign csr_io_rocc_autl_acquire_valid = GEN_257;
  assign csr_io_rocc_autl_acquire_bits_addr_block = GEN_258;
  assign csr_io_rocc_autl_acquire_bits_client_xact_id = GEN_259;
  assign csr_io_rocc_autl_acquire_bits_addr_beat = GEN_260;
  assign csr_io_rocc_autl_acquire_bits_is_builtin_type = GEN_261;
  assign csr_io_rocc_autl_acquire_bits_a_type = GEN_262;
  assign csr_io_rocc_autl_acquire_bits_union = GEN_263;
  assign csr_io_rocc_autl_acquire_bits_data = GEN_264;
  assign csr_io_rocc_autl_grant_ready = GEN_265;
  assign csr_io_rocc_fpu_req_valid = GEN_266;
  assign csr_io_rocc_fpu_req_bits_cmd = GEN_267;
  assign csr_io_rocc_fpu_req_bits_ldst = GEN_268;
  assign csr_io_rocc_fpu_req_bits_wen = GEN_269;
  assign csr_io_rocc_fpu_req_bits_ren1 = GEN_270;
  assign csr_io_rocc_fpu_req_bits_ren2 = GEN_271;
  assign csr_io_rocc_fpu_req_bits_ren3 = GEN_272;
  assign csr_io_rocc_fpu_req_bits_swap12 = GEN_273;
  assign csr_io_rocc_fpu_req_bits_swap23 = GEN_274;
  assign csr_io_rocc_fpu_req_bits_single = GEN_275;
  assign csr_io_rocc_fpu_req_bits_fromint = GEN_276;
  assign csr_io_rocc_fpu_req_bits_toint = GEN_277;
  assign csr_io_rocc_fpu_req_bits_fastpipe = GEN_278;
  assign csr_io_rocc_fpu_req_bits_fma = GEN_279;
  assign csr_io_rocc_fpu_req_bits_div = GEN_280;
  assign csr_io_rocc_fpu_req_bits_sqrt = GEN_281;
  assign csr_io_rocc_fpu_req_bits_round = GEN_282;
  assign csr_io_rocc_fpu_req_bits_wflags = GEN_283;
  assign csr_io_rocc_fpu_req_bits_rm = GEN_284;
  assign csr_io_rocc_fpu_req_bits_typ = GEN_285;
  assign csr_io_rocc_fpu_req_bits_in1 = GEN_286;
  assign csr_io_rocc_fpu_req_bits_in2 = GEN_287;
  assign csr_io_rocc_fpu_req_bits_in3 = GEN_288;
  assign csr_io_rocc_fpu_resp_ready = GEN_289;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign T_7207 = id_ctrl_csr == 3'h2;
  assign T_7208 = id_ctrl_csr == 3'h3;
  assign T_7209 = T_7207 | T_7208;
  assign id_csr_ren = T_7209 & T_7188;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_csr_addr = io_imem_resp_bits_data_0[31:20];
  assign T_7213 = id_csr_ren == 1'h0;
  assign T_7214 = id_csr_en & T_7213;
  assign T_7268 = id_csr_addr & 12'h46;
  assign T_7270 = T_7268 == 12'h40;
  assign T_7272 = id_csr_addr & 12'h644;
  assign T_7274 = T_7272 == 12'h240;
  assign T_7277 = T_7270 | T_7274;
  assign T_7280 = T_7277 == 1'h0;
  assign T_7281 = T_7214 & T_7280;
  assign id_csr_flush = id_system_insn | T_7281;
  assign T_7283 = id_ctrl_legal == 1'h0;
  assign GEN_173 = {{1'd0}, 1'h0};
  assign T_7285 = csr_io_status_fs != GEN_173;
  assign T_7287 = T_7285 == 1'h0;
  assign T_7288 = id_ctrl_fp & T_7287;
  assign T_7289 = T_7283 | T_7288;
  assign T_7291 = csr_io_status_xs != GEN_173;
  assign T_7293 = T_7291 == 1'h0;
  assign T_7294 = id_ctrl_rocc & T_7293;
  assign id_illegal_insn = T_7289 | T_7294;
  assign id_amo_aq = io_imem_resp_bits_data_0[26];
  assign id_amo_rl = io_imem_resp_bits_data_0[25];
  assign T_7295 = id_ctrl_amo & id_amo_rl;
  assign id_fence_next = id_ctrl_fence | T_7295;
  assign T_7297 = io_dmem_ordered == 1'h0;
  assign id_mem_busy = T_7297 | io_dmem_req_valid;
  assign T_7303 = wb_reg_valid & wb_ctrl_rocc;
  assign T_7305 = id_reg_fence & id_mem_busy;
  assign T_7306 = id_fence_next | T_7305;
  assign T_7308 = id_ctrl_amo & id_amo_aq;
  assign T_7309 = T_7308 | id_ctrl_fence_i;
  assign T_7310 = id_ctrl_mem | id_ctrl_rocc;
  assign T_7311 = id_reg_fence & T_7310;
  assign T_7312 = T_7309 | T_7311;
  assign T_7313 = T_7312 | id_csr_en;
  assign T_7314 = id_mem_busy & T_7313;
  assign bpu_clk = clk;
  assign bpu_reset = reset;
  assign bpu_io_status_debug = csr_io_status_debug;
  assign bpu_io_status_prv = csr_io_status_prv;
  assign bpu_io_status_sd = csr_io_status_sd;
  assign bpu_io_status_zero3 = csr_io_status_zero3;
  assign bpu_io_status_sd_rv32 = csr_io_status_sd_rv32;
  assign bpu_io_status_zero2 = csr_io_status_zero2;
  assign bpu_io_status_vm = csr_io_status_vm;
  assign bpu_io_status_zero1 = csr_io_status_zero1;
  assign bpu_io_status_pum = csr_io_status_pum;
  assign bpu_io_status_mprv = csr_io_status_mprv;
  assign bpu_io_status_xs = csr_io_status_xs;
  assign bpu_io_status_fs = csr_io_status_fs;
  assign bpu_io_status_mpp = csr_io_status_mpp;
  assign bpu_io_status_hpp = csr_io_status_hpp;
  assign bpu_io_status_spp = csr_io_status_spp;
  assign bpu_io_status_mpie = csr_io_status_mpie;
  assign bpu_io_status_hpie = csr_io_status_hpie;
  assign bpu_io_status_spie = csr_io_status_spie;
  assign bpu_io_status_upie = csr_io_status_upie;
  assign bpu_io_status_mie = csr_io_status_mie;
  assign bpu_io_status_hie = csr_io_status_hie;
  assign bpu_io_status_sie = csr_io_status_sie;
  assign bpu_io_status_uie = csr_io_status_uie;
  assign bpu_io_bp_0_control_tdrtype = csr_io_bp_0_control_tdrtype;
  assign bpu_io_bp_0_control_bpamaskmax = csr_io_bp_0_control_bpamaskmax;
  assign bpu_io_bp_0_control_reserved = csr_io_bp_0_control_reserved;
  assign bpu_io_bp_0_control_bpaction = csr_io_bp_0_control_bpaction;
  assign bpu_io_bp_0_control_bpmatch = csr_io_bp_0_control_bpmatch;
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m;
  assign bpu_io_bp_0_control_h = csr_io_bp_0_control_h;
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s;
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u;
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r;
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w;
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x;
  assign bpu_io_bp_0_address = csr_io_bp_0_address;
  assign bpu_io_pc = io_imem_resp_bits_pc[38:0];
  assign bpu_io_ea = mem_reg_wdata[38:0];
  assign T_7318 = csr_io_interrupt | bpu_io_xcpt_if;
  assign T_7319 = T_7318 | io_imem_resp_bits_xcpt_if;
  assign id_xcpt = T_7319 | id_illegal_insn;
  assign T_7320 = io_imem_resp_bits_xcpt_if ? {{1'd0}, 1'h1} : 2'h2;
  assign T_7321 = bpu_io_xcpt_if ? 2'h3 : T_7320;
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : {{62'd0}, T_7321};
  assign ex_waddr = ex_reg_inst[11:7];
  assign mem_waddr = mem_reg_inst[11:7];
  assign wb_waddr = wb_reg_inst[11:7];
  assign T_7325 = ex_reg_valid & ex_ctrl_wxd;
  assign T_7326 = mem_reg_valid & mem_ctrl_wxd;
  assign T_7328 = mem_ctrl_mem == 1'h0;
  assign T_7329 = T_7326 & T_7328;
  assign T_7331 = GEN_170 == id_raddr1;
  assign T_7333 = ex_waddr == id_raddr1;
  assign T_7334 = T_7325 & T_7333;
  assign T_7335 = mem_waddr == id_raddr1;
  assign T_7336 = T_7329 & T_7335;
  assign T_7338 = T_7326 & T_7335;
  assign T_7339 = GEN_170 == id_raddr2;
  assign T_7341 = ex_waddr == id_raddr2;
  assign T_7342 = T_7325 & T_7341;
  assign T_7343 = mem_waddr == id_raddr2;
  assign T_7344 = T_7329 & T_7343;
  assign T_7346 = T_7326 & T_7343;
  assign bypass_mux_0 = {{63'd0}, 1'h0};
  assign bypass_mux_1 = mem_reg_wdata;
  assign bypass_mux_2 = wb_reg_wdata;
  assign bypass_mux_3 = io_dmem_resp_bits_data_word_bypass;
  assign T_7374 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0};
  assign GEN_0 = GEN_4;
  assign GEN_177 = {{1'd0}, 1'h1};
  assign GEN_2 = GEN_177 == ex_reg_rs_lsb_0 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_3 = 2'h2 == ex_reg_rs_lsb_0 ? bypass_mux_2 : GEN_2;
  assign GEN_4 = 2'h3 == ex_reg_rs_lsb_0 ? bypass_mux_3 : GEN_3;
  assign T_7375 = ex_reg_rs_bypass_0 ? GEN_0 : T_7374;
  assign T_7376 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1};
  assign GEN_1 = GEN_7;
  assign GEN_5 = GEN_177 == ex_reg_rs_lsb_1 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_6 = 2'h2 == ex_reg_rs_lsb_1 ? bypass_mux_2 : GEN_5;
  assign GEN_7 = 2'h3 == ex_reg_rs_lsb_1 ? bypass_mux_3 : GEN_6;
  assign T_7377 = ex_reg_rs_bypass_1 ? GEN_1 : T_7376;
  assign T_7378 = ex_ctrl_sel_imm == 3'h5;
  assign T_7380 = ex_reg_inst[31];
  assign T_7381 = $signed(T_7380);
  assign T_7382 = T_7378 ? $signed($signed(1'h0)) : $signed(T_7381);
  assign T_7383 = ex_ctrl_sel_imm == 3'h2;
  assign T_7384 = ex_reg_inst[30:20];
  assign T_7385 = $signed(T_7384);
  assign T_7386 = T_7383 ? $signed(T_7385) : $signed({11{T_7382}});
  assign T_7387 = ex_ctrl_sel_imm != 3'h2;
  assign T_7388 = ex_ctrl_sel_imm != 3'h3;
  assign T_7389 = T_7387 & T_7388;
  assign T_7390 = ex_reg_inst[19:12];
  assign T_7391 = $signed(T_7390);
  assign T_7392 = T_7389 ? $signed({8{T_7382}}) : $signed(T_7391);
  assign T_7395 = T_7383 | T_7378;
  assign T_7397 = ex_ctrl_sel_imm == 3'h3;
  assign T_7398 = ex_reg_inst[20];
  assign T_7399 = $signed(T_7398);
  assign T_7400 = ex_ctrl_sel_imm == 3'h1;
  assign T_7401 = ex_reg_inst[7];
  assign T_7402 = $signed(T_7401);
  assign T_7403 = T_7400 ? $signed(T_7402) : $signed(T_7382);
  assign T_7404 = T_7397 ? $signed(T_7399) : $signed(T_7403);
  assign T_7405 = T_7395 ? $signed($signed(1'h0)) : $signed(T_7404);
  assign T_7410 = ex_reg_inst[30:25];
  assign T_7411 = T_7395 ? {{5'd0}, 1'h0} : T_7410;
  assign T_7414 = ex_ctrl_sel_imm == 3'h0;
  assign T_7416 = T_7414 | T_7400;
  assign T_7417 = ex_reg_inst[11:8];
  assign T_7419 = ex_reg_inst[19:16];
  assign T_7420 = ex_reg_inst[24:21];
  assign T_7421 = T_7378 ? T_7419 : T_7420;
  assign T_7422 = T_7416 ? T_7417 : T_7421;
  assign T_7423 = T_7383 ? {{3'd0}, 1'h0} : T_7422;
  assign T_7426 = ex_ctrl_sel_imm == 3'h4;
  assign T_7429 = ex_reg_inst[15];
  assign T_7432 = T_7378 ? T_7429 : 1'h0;
  assign T_7434 = T_7426 ? T_7398 : T_7432;
  assign T_7436 = T_7414 ? T_7401 : T_7434;
  assign T_7437 = {T_7411,T_7423};
  assign T_7438 = {T_7437,T_7436};
  assign T_7439 = $unsigned(T_7405);
  assign T_7440 = $unsigned(T_7392);
  assign T_7441 = {T_7440,T_7439};
  assign T_7442 = $unsigned(T_7386);
  assign T_7443 = $unsigned(T_7382);
  assign T_7444 = {T_7443,T_7442};
  assign T_7445 = {T_7444,T_7441};
  assign T_7446 = {T_7445,T_7438};
  assign ex_imm = $signed(T_7446);
  assign T_7448 = $signed(T_7375);
  assign T_7449 = $signed(ex_reg_pc);
  assign T_7450 = 2'h2 == ex_ctrl_sel_alu1;
  assign GEN_179 = $signed(1'h0);
  assign T_7451 = T_7450 ? $signed(T_7449) : $signed({40{GEN_179}});
  assign T_7452 = 2'h1 == ex_ctrl_sel_alu1;
  assign ex_op1 = T_7452 ? $signed(T_7448) : $signed({{24{T_7451[39]}},T_7451});
  assign T_7454 = $signed(T_7377);
  assign T_7456 = 2'h1 == ex_ctrl_sel_alu2;
  assign T_7457 = T_7456 ? $signed($signed(4'h4)) : $signed({4{GEN_179}});
  assign T_7458 = 2'h3 == ex_ctrl_sel_alu2;
  assign T_7459 = T_7458 ? $signed(ex_imm) : $signed({{28{T_7457[3]}},T_7457});
  assign T_7460 = 2'h2 == ex_ctrl_sel_alu2;
  assign ex_op2 = T_7460 ? $signed(T_7454) : $signed({{32{T_7459[31]}},T_7459});
  assign alu_clk = clk;
  assign alu_reset = reset;
  assign alu_io_dw = ex_ctrl_alu_dw;
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign alu_io_in2 = T_7461;
  assign alu_io_in1 = T_7462;
  assign T_7461 = $unsigned(ex_op2);
  assign T_7462 = $unsigned(ex_op1);
  assign div_clk = clk;
  assign div_reset = reset;
  assign div_io_req_valid = T_7463;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_dw = ex_ctrl_alu_dw;
  assign div_io_req_bits_in1 = T_7375;
  assign div_io_req_bits_in2 = T_7377;
  assign div_io_req_bits_tag = ex_waddr;
  assign div_io_kill = T_7800;
  assign div_io_resp_ready = GEN_149;
  assign T_7463 = ex_reg_valid & ex_ctrl_div;
  assign T_7465 = ctrl_killd == 1'h0;
  assign T_7468 = T_7465 & id_xcpt;
  assign T_7470 = take_pc_mem_wb == 1'h0;
  assign T_7471 = csr_io_interrupt & T_7470;
  assign T_7472 = T_7471 & io_imem_resp_valid;
  assign GEN_8 = id_xcpt ? id_cause : ex_reg_cause;
  assign GEN_9 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign GEN_10 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_mask : ex_reg_btb_resp_mask;
  assign GEN_11 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bridx : ex_reg_btb_resp_bridx;
  assign GEN_12 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign GEN_13 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign GEN_14 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign GEN_15 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T_7475 = id_ctrl_fence_i | id_csr_flush;
  assign T_7476 = T_7475 | csr_io_singleStep;
  assign T_7477 = id_ctrl_jalr & csr_io_status_debug;
  assign GEN_16 = T_7477 ? 1'h1 : T_7476;
  assign GEN_17 = T_7477 ? 1'h1 : id_ctrl_fence_i;
  assign T_7480 = T_7331 | T_7334;
  assign T_7481 = T_7480 | T_7336;
  assign T_7482 = T_7481 | T_7338;
  assign T_7487 = T_7336 ? 2'h2 : 2'h3;
  assign T_7488 = T_7334 ? {{1'd0}, 1'h1} : T_7487;
  assign T_7489 = T_7331 ? {{1'd0}, 1'h0} : T_7488;
  assign T_7491 = T_7482 == 1'h0;
  assign T_7492 = id_ctrl_rxs1 & T_7491;
  assign T_7493 = T_7185[1:0];
  assign T_7494 = T_7185[63:2];
  assign GEN_18 = T_7492 ? T_7493 : T_7489;
  assign GEN_19 = T_7492 ? T_7494 : ex_reg_rs_msb_0;
  assign T_7495 = T_7339 | T_7342;
  assign T_7496 = T_7495 | T_7344;
  assign T_7497 = T_7496 | T_7346;
  assign T_7502 = T_7344 ? 2'h2 : 2'h3;
  assign T_7503 = T_7342 ? {{1'd0}, 1'h1} : T_7502;
  assign T_7504 = T_7339 ? {{1'd0}, 1'h0} : T_7503;
  assign T_7506 = T_7497 == 1'h0;
  assign T_7507 = id_ctrl_rxs2 & T_7506;
  assign T_7508 = T_7196[1:0];
  assign T_7509 = T_7196[63:2];
  assign GEN_20 = T_7507 ? T_7508 : T_7504;
  assign GEN_21 = T_7507 ? T_7509 : ex_reg_rs_msb_1;
  assign GEN_22 = T_7465 ? id_ctrl_legal : ex_ctrl_legal;
  assign GEN_23 = T_7465 ? id_ctrl_fp : ex_ctrl_fp;
  assign GEN_24 = T_7465 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign GEN_25 = T_7465 ? id_ctrl_branch : ex_ctrl_branch;
  assign GEN_26 = T_7465 ? id_ctrl_jal : ex_ctrl_jal;
  assign GEN_27 = T_7465 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign GEN_28 = T_7465 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign GEN_29 = T_7465 ? id_ctrl_rxs1 : ex_ctrl_rxs1;
  assign GEN_30 = T_7465 ? id_ctrl_sel_alu2 : ex_ctrl_sel_alu2;
  assign GEN_31 = T_7465 ? id_ctrl_sel_alu1 : ex_ctrl_sel_alu1;
  assign GEN_32 = T_7465 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign GEN_33 = T_7465 ? id_ctrl_alu_dw : ex_ctrl_alu_dw;
  assign GEN_34 = T_7465 ? id_ctrl_alu_fn : ex_ctrl_alu_fn;
  assign GEN_35 = T_7465 ? id_ctrl_mem : ex_ctrl_mem;
  assign GEN_36 = T_7465 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign GEN_37 = T_7465 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign GEN_38 = T_7465 ? id_ctrl_rfs1 : ex_ctrl_rfs1;
  assign GEN_39 = T_7465 ? id_ctrl_rfs2 : ex_ctrl_rfs2;
  assign GEN_40 = T_7465 ? id_ctrl_rfs3 : ex_ctrl_rfs3;
  assign GEN_41 = T_7465 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign GEN_42 = T_7465 ? id_ctrl_div : ex_ctrl_div;
  assign GEN_43 = T_7465 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign GEN_44 = T_7465 ? id_csr : ex_ctrl_csr;
  assign GEN_45 = T_7465 ? GEN_17 : ex_ctrl_fence_i;
  assign GEN_46 = T_7465 ? id_ctrl_fence : ex_ctrl_fence;
  assign GEN_47 = T_7465 ? id_ctrl_amo : ex_ctrl_amo;
  assign GEN_48 = T_7465 ? io_imem_btb_resp_valid : ex_reg_btb_hit;
  assign GEN_49 = T_7465 ? GEN_9 : ex_reg_btb_resp_taken;
  assign GEN_50 = T_7465 ? GEN_10 : ex_reg_btb_resp_mask;
  assign GEN_51 = T_7465 ? GEN_11 : ex_reg_btb_resp_bridx;
  assign GEN_52 = T_7465 ? GEN_12 : ex_reg_btb_resp_target;
  assign GEN_53 = T_7465 ? GEN_13 : ex_reg_btb_resp_entry;
  assign GEN_54 = T_7465 ? GEN_14 : ex_reg_btb_resp_bht_history;
  assign GEN_55 = T_7465 ? GEN_15 : ex_reg_btb_resp_bht_value;
  assign GEN_56 = T_7465 ? GEN_16 : ex_reg_flush_pipe;
  assign GEN_57 = T_7465 ? id_load_use : ex_reg_load_use;
  assign GEN_58 = T_7465 ? T_7482 : ex_reg_rs_bypass_0;
  assign GEN_59 = T_7465 ? GEN_18 : ex_reg_rs_lsb_0;
  assign GEN_60 = T_7465 ? GEN_19 : ex_reg_rs_msb_0;
  assign GEN_61 = T_7465 ? T_7497 : ex_reg_rs_bypass_1;
  assign GEN_62 = T_7465 ? GEN_20 : ex_reg_rs_lsb_1;
  assign GEN_63 = T_7465 ? GEN_21 : ex_reg_rs_msb_1;
  assign T_7512 = T_7465 | csr_io_interrupt;
  assign GEN_64 = T_7512 ? io_imem_resp_bits_data_0 : ex_reg_inst;
  assign GEN_65 = T_7512 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign ex_pc_valid = ex_reg_valid | ex_reg_xcpt_interrupt;
  assign T_7514 = io_dmem_resp_valid == 1'h0;
  assign wb_dcache_miss = wb_ctrl_mem & T_7514;
  assign T_7516 = io_dmem_req_ready == 1'h0;
  assign T_7517 = ex_ctrl_mem & T_7516;
  assign T_7519 = div_io_req_ready == 1'h0;
  assign T_7520 = ex_ctrl_div & T_7519;
  assign replay_ex_structural = T_7517 | T_7520;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T_7521 = replay_ex_structural | replay_ex_load_use;
  assign replay_ex = ex_reg_valid & T_7521;
  assign T_7522 = take_pc_mem_wb | replay_ex;
  assign T_7524 = ex_reg_valid == 1'h0;
  assign ctrl_killx = T_7522 | T_7524;
  assign T_7525 = ex_ctrl_mem_cmd == 5'h7;
  assign T_7531_0 = 3'h0;
  assign T_7531_1 = 3'h4;
  assign T_7531_2 = 3'h1;
  assign T_7531_3 = 3'h5;
  assign T_7533 = T_7531_0 == ex_ctrl_mem_type;
  assign T_7534 = T_7531_1 == ex_ctrl_mem_type;
  assign T_7535 = T_7531_2 == ex_ctrl_mem_type;
  assign T_7536 = T_7531_3 == ex_ctrl_mem_type;
  assign T_7539 = T_7533 | T_7534;
  assign T_7540 = T_7539 | T_7535;
  assign T_7541 = T_7540 | T_7536;
  assign ex_slow_bypass = T_7525 | T_7541;
  assign T_7542 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T_7543 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign ex_xcpt = T_7542 | T_7543;
  assign ex_cause = T_7542 ? ex_reg_cause : {{62'd0}, 2'h2};
  assign mem_br_taken = mem_reg_wdata[0];
  assign T_7545 = $signed(mem_reg_pc);
  assign T_7546 = mem_ctrl_branch & mem_br_taken;
  assign T_7549 = mem_reg_inst[31];
  assign T_7550 = $signed(T_7549);
  assign T_7551 = 1'h0 ? $signed($signed(1'h0)) : $signed(T_7550);
  assign T_7553 = mem_reg_inst[30:20];
  assign T_7554 = $signed(T_7553);
  assign T_7555 = 1'h0 ? $signed(T_7554) : $signed({11{T_7551}});
  assign T_7559 = mem_reg_inst[19:12];
  assign T_7560 = $signed(T_7559);
  assign T_7561 = 1'h1 ? $signed({8{T_7551}}) : $signed(T_7560);
  assign T_7567 = mem_reg_inst[20];
  assign T_7568 = $signed(T_7567);
  assign T_7570 = mem_reg_inst[7];
  assign T_7571 = $signed(T_7570);
  assign T_7572 = 1'h1 ? $signed(T_7571) : $signed(T_7551);
  assign T_7573 = 1'h0 ? $signed(T_7568) : $signed(T_7572);
  assign T_7574 = 1'h0 ? $signed($signed(1'h0)) : $signed(T_7573);
  assign T_7579 = mem_reg_inst[30:25];
  assign T_7586 = mem_reg_inst[11:8];
  assign T_7589 = mem_reg_inst[24:21];
  assign T_7606 = {T_7579,T_7586};
  assign T_7607 = {T_7606,1'h0};
  assign T_7608 = $unsigned(T_7574);
  assign T_7609 = $unsigned(T_7561);
  assign T_7610 = {T_7609,T_7608};
  assign T_7611 = $unsigned(T_7555);
  assign T_7612 = $unsigned(T_7551);
  assign T_7613 = {T_7612,T_7611};
  assign T_7614 = {T_7613,T_7610};
  assign T_7615 = {T_7614,T_7607};
  assign T_7616 = $signed(T_7615);
  assign T_7631 = 1'h0 ? $signed({8{T_7551}}) : $signed(T_7560);
  assign T_7642 = 1'h0 ? $signed(T_7571) : $signed(T_7551);
  assign T_7643 = 1'h1 ? $signed(T_7568) : $signed(T_7642);
  assign T_7644 = 1'h0 ? $signed($signed(1'h0)) : $signed(T_7643);
  assign T_7676 = {T_7579,T_7589};
  assign T_7677 = {T_7676,1'h0};
  assign T_7678 = $unsigned(T_7644);
  assign T_7679 = $unsigned(T_7631);
  assign T_7680 = {T_7679,T_7678};
  assign T_7684 = {T_7613,T_7680};
  assign T_7685 = {T_7684,T_7677};
  assign T_7686 = $signed(T_7685);
  assign GEN_181 = $signed(4'h4);
  assign T_7688 = mem_ctrl_jal ? $signed(T_7686) : $signed({{28{GEN_181[3]}},GEN_181});
  assign T_7689 = T_7546 ? $signed(T_7616) : $signed(T_7688);
  assign GEN_182 = {{8{T_7689[31]}},T_7689};
  assign T_7690 = $signed(T_7545) + $signed(GEN_182);
  assign T_7691 = T_7690[39:0];
  assign mem_br_target = $signed(T_7691);
  assign T_7692 = $signed(mem_reg_wdata);
  assign T_7693 = mem_ctrl_jalr ? $signed({{24{mem_br_target[39]}},mem_br_target}) : $signed(T_7692);
  assign mem_int_wdata = $unsigned(T_7693);
  assign T_7694 = mem_reg_wdata[63:38];
  assign T_7695 = mem_reg_wdata[39:38];
  assign T_7696 = $signed(T_7695);
  assign GEN_183 = {{25'd0}, 1'h0};
  assign T_7698 = T_7694 == GEN_183;
  assign GEN_184 = {{25'd0}, 1'h1};
  assign T_7700 = T_7694 == GEN_184;
  assign T_7701 = T_7698 | T_7700;
  assign GEN_186 = {2{GEN_179}};
  assign T_7703 = $signed(T_7696) != $signed(GEN_186);
  assign T_7704 = $signed(T_7694);
  assign GEN_187 = $signed(1'h1);
  assign GEN_188 = {26{GEN_187}};
  assign T_7706 = $signed(T_7704) == $signed(GEN_188);
  assign GEN_189 = $signed(2'h2);
  assign GEN_190 = {{24{GEN_189[1]}},GEN_189};
  assign T_7709 = $signed(T_7704) == $signed(GEN_190);
  assign T_7710 = T_7706 | T_7709;
  assign GEN_192 = {2{GEN_187}};
  assign T_7712 = $signed(T_7696) == $signed(GEN_192);
  assign T_7713 = T_7696[0];
  assign T_7714 = T_7710 ? T_7712 : T_7713;
  assign T_7715 = T_7701 ? T_7703 : T_7714;
  assign T_7716 = mem_reg_wdata[38:0];
  assign T_7717 = {T_7715,T_7716};
  assign T_7718 = $signed(T_7717);
  assign T_7719 = mem_ctrl_jalr ? $signed(T_7718) : $signed(mem_br_target);
  assign GEN_194 = {{38{GEN_189[1]}},GEN_189};
  assign T_7721 = $signed(T_7719) & $signed(GEN_194);
  assign T_7722 = $signed(T_7721);
  assign mem_npc = $unsigned(T_7722);
  assign T_7723 = mem_npc != ex_reg_pc;
  assign T_7724 = mem_npc != io_imem_resp_bits_pc;
  assign T_7726 = io_imem_resp_valid ? T_7724 : 1'h1;
  assign mem_wrong_npc = ex_pc_valid ? T_7723 : T_7726;
  assign mem_npc_misaligned = mem_npc[1];
  assign T_7729 = T_7546 | mem_ctrl_jalr;
  assign mem_cfi_taken = T_7729 | mem_ctrl_jal;
  assign T_7730 = mem_wrong_npc | mem_reg_flush_pipe;
  assign want_take_pc_mem = mem_reg_valid & T_7730;
  assign T_7732 = mem_npc_misaligned == 1'h0;
  assign T_7733 = want_take_pc_mem & T_7732;
  assign T_7735 = ctrl_killx == 1'h0;
  assign T_7738 = T_7470 & replay_ex;
  assign T_7741 = T_7735 & ex_xcpt;
  assign T_7744 = T_7470 & ex_reg_xcpt_interrupt;
  assign GEN_66 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign T_7745 = ex_ctrl_mem_cmd == 5'h0;
  assign T_7746 = ex_ctrl_mem_cmd == 5'h6;
  assign T_7747 = T_7745 | T_7746;
  assign T_7749 = T_7747 | T_7525;
  assign T_7750 = ex_ctrl_mem_cmd[3];
  assign T_7751 = ex_ctrl_mem_cmd == 5'h4;
  assign T_7752 = T_7750 | T_7751;
  assign T_7753 = T_7749 | T_7752;
  assign T_7754 = ex_ctrl_mem & T_7753;
  assign T_7755 = ex_ctrl_mem_cmd == 5'h1;
  assign T_7757 = T_7755 | T_7525;
  assign T_7761 = T_7757 | T_7752;
  assign T_7762 = ex_ctrl_mem & T_7761;
  assign GEN_67 = ex_reg_btb_hit ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign GEN_68 = ex_reg_btb_hit ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign GEN_69 = ex_reg_btb_hit ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign GEN_70 = ex_reg_btb_hit ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign GEN_71 = ex_reg_btb_hit ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign GEN_72 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign GEN_73 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T_7763 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T_7764 = ex_ctrl_rxs2 & T_7763;
  assign GEN_74 = T_7764 ? T_7377 : mem_reg_rs2;
  assign GEN_75 = ex_pc_valid ? ex_ctrl_legal : mem_ctrl_legal;
  assign GEN_76 = ex_pc_valid ? ex_ctrl_fp : mem_ctrl_fp;
  assign GEN_77 = ex_pc_valid ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign GEN_78 = ex_pc_valid ? ex_ctrl_branch : mem_ctrl_branch;
  assign GEN_79 = ex_pc_valid ? ex_ctrl_jal : mem_ctrl_jal;
  assign GEN_80 = ex_pc_valid ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign GEN_81 = ex_pc_valid ? ex_ctrl_rxs2 : mem_ctrl_rxs2;
  assign GEN_82 = ex_pc_valid ? ex_ctrl_rxs1 : mem_ctrl_rxs1;
  assign GEN_83 = ex_pc_valid ? ex_ctrl_sel_alu2 : mem_ctrl_sel_alu2;
  assign GEN_84 = ex_pc_valid ? ex_ctrl_sel_alu1 : mem_ctrl_sel_alu1;
  assign GEN_85 = ex_pc_valid ? ex_ctrl_sel_imm : mem_ctrl_sel_imm;
  assign GEN_86 = ex_pc_valid ? ex_ctrl_alu_dw : mem_ctrl_alu_dw;
  assign GEN_87 = ex_pc_valid ? ex_ctrl_alu_fn : mem_ctrl_alu_fn;
  assign GEN_88 = ex_pc_valid ? ex_ctrl_mem : mem_ctrl_mem;
  assign GEN_89 = ex_pc_valid ? ex_ctrl_mem_cmd : mem_ctrl_mem_cmd;
  assign GEN_90 = ex_pc_valid ? ex_ctrl_mem_type : mem_ctrl_mem_type;
  assign GEN_91 = ex_pc_valid ? ex_ctrl_rfs1 : mem_ctrl_rfs1;
  assign GEN_92 = ex_pc_valid ? ex_ctrl_rfs2 : mem_ctrl_rfs2;
  assign GEN_93 = ex_pc_valid ? ex_ctrl_rfs3 : mem_ctrl_rfs3;
  assign GEN_94 = ex_pc_valid ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign GEN_95 = ex_pc_valid ? ex_ctrl_div : mem_ctrl_div;
  assign GEN_96 = ex_pc_valid ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign GEN_97 = ex_pc_valid ? ex_ctrl_csr : mem_ctrl_csr;
  assign GEN_98 = ex_pc_valid ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign GEN_99 = ex_pc_valid ? ex_ctrl_fence : mem_ctrl_fence;
  assign GEN_100 = ex_pc_valid ? ex_ctrl_amo : mem_ctrl_amo;
  assign GEN_101 = ex_pc_valid ? T_7754 : mem_reg_load;
  assign GEN_102 = ex_pc_valid ? T_7762 : mem_reg_store;
  assign GEN_103 = ex_pc_valid ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign GEN_104 = ex_pc_valid ? GEN_67 : mem_reg_btb_resp_taken;
  assign GEN_105 = ex_pc_valid ? GEN_68 : mem_reg_btb_resp_mask;
  assign GEN_106 = ex_pc_valid ? GEN_69 : mem_reg_btb_resp_bridx;
  assign GEN_107 = ex_pc_valid ? GEN_70 : mem_reg_btb_resp_target;
  assign GEN_108 = ex_pc_valid ? GEN_71 : mem_reg_btb_resp_entry;
  assign GEN_109 = ex_pc_valid ? GEN_72 : mem_reg_btb_resp_bht_history;
  assign GEN_110 = ex_pc_valid ? GEN_73 : mem_reg_btb_resp_bht_value;
  assign GEN_111 = ex_pc_valid ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign GEN_112 = ex_pc_valid ? ex_slow_bypass : mem_reg_slow_bypass;
  assign GEN_113 = ex_pc_valid ? ex_reg_inst : mem_reg_inst;
  assign GEN_114 = ex_pc_valid ? ex_reg_pc : mem_reg_pc;
  assign GEN_115 = ex_pc_valid ? alu_io_out : mem_reg_wdata;
  assign GEN_116 = ex_pc_valid ? GEN_74 : mem_reg_rs2;
  assign T_7765 = mem_reg_load & bpu_io_xcpt_ld;
  assign T_7767 = mem_reg_store & bpu_io_xcpt_st;
  assign T_7769 = want_take_pc_mem & mem_npc_misaligned;
  assign T_7771 = mem_ctrl_mem & io_dmem_xcpt_ma_st;
  assign T_7773 = mem_ctrl_mem & io_dmem_xcpt_ma_ld;
  assign T_7775 = mem_ctrl_mem & io_dmem_xcpt_pf_st;
  assign T_7777 = mem_ctrl_mem & io_dmem_xcpt_pf_ld;
  assign T_7779 = T_7765 | T_7767;
  assign T_7780 = T_7779 | T_7769;
  assign T_7781 = T_7780 | T_7771;
  assign T_7782 = T_7781 | T_7773;
  assign T_7783 = T_7782 | T_7775;
  assign mem_new_xcpt = T_7783 | T_7777;
  assign T_7784 = T_7775 ? 3'h7 : 3'h5;
  assign T_7785 = T_7773 ? 3'h4 : T_7784;
  assign T_7786 = T_7771 ? 3'h6 : T_7785;
  assign T_7787 = T_7769 ? {{2'd0}, 1'h0} : T_7786;
  assign T_7788 = T_7767 ? {{1'd0}, 2'h3} : T_7787;
  assign mem_new_cause = T_7765 ? {{1'd0}, 2'h3} : T_7788;
  assign T_7789 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T_7790 = mem_reg_valid & mem_new_xcpt;
  assign mem_xcpt = T_7789 | T_7790;
  assign mem_cause = T_7789 ? mem_reg_cause : {{61'd0}, mem_new_cause};
  assign dcache_kill_mem = T_7326 & io_dmem_replay_next;
  assign T_7792 = mem_reg_valid & mem_ctrl_fp;
  assign fpu_kill_mem = T_7792 & io_fpu_nack_mem;
  assign T_7793 = dcache_kill_mem | mem_reg_replay;
  assign replay_mem = T_7793 | fpu_kill_mem;
  assign T_7794 = dcache_kill_mem | take_pc_wb;
  assign T_7795 = T_7794 | mem_reg_xcpt;
  assign T_7797 = mem_reg_valid == 1'h0;
  assign killm_common = T_7795 | T_7797;
  assign T_7798 = div_io_req_ready & div_io_req_valid;
  assign T_7800 = killm_common & T_7799;
  assign T_7801 = killm_common | mem_xcpt;
  assign ctrl_killm = T_7801 | fpu_kill_mem;
  assign T_7803 = ctrl_killm == 1'h0;
  assign T_7805 = take_pc_wb == 1'h0;
  assign T_7806 = replay_mem & T_7805;
  assign T_7809 = mem_xcpt & T_7805;
  assign T_7813 = T_7789 == 1'h0;
  assign T_7814 = T_7790 & T_7813;
  assign GEN_117 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign T_7815 = mem_reg_valid | mem_reg_replay;
  assign T_7816 = T_7815 | mem_reg_xcpt_interrupt;
  assign T_7817 = mem_ctrl_fp & mem_ctrl_wxd;
  assign T_7818 = T_7817 ? io_fpu_toint_data : mem_int_wdata;
  assign GEN_118 = mem_ctrl_rocc ? mem_reg_rs2 : wb_reg_rs2;
  assign GEN_119 = T_7816 ? mem_ctrl_legal : wb_ctrl_legal;
  assign GEN_120 = T_7816 ? mem_ctrl_fp : wb_ctrl_fp;
  assign GEN_121 = T_7816 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign GEN_122 = T_7816 ? mem_ctrl_branch : wb_ctrl_branch;
  assign GEN_123 = T_7816 ? mem_ctrl_jal : wb_ctrl_jal;
  assign GEN_124 = T_7816 ? mem_ctrl_jalr : wb_ctrl_jalr;
  assign GEN_125 = T_7816 ? mem_ctrl_rxs2 : wb_ctrl_rxs2;
  assign GEN_126 = T_7816 ? mem_ctrl_rxs1 : wb_ctrl_rxs1;
  assign GEN_127 = T_7816 ? mem_ctrl_sel_alu2 : wb_ctrl_sel_alu2;
  assign GEN_128 = T_7816 ? mem_ctrl_sel_alu1 : wb_ctrl_sel_alu1;
  assign GEN_129 = T_7816 ? mem_ctrl_sel_imm : wb_ctrl_sel_imm;
  assign GEN_130 = T_7816 ? mem_ctrl_alu_dw : wb_ctrl_alu_dw;
  assign GEN_131 = T_7816 ? mem_ctrl_alu_fn : wb_ctrl_alu_fn;
  assign GEN_132 = T_7816 ? mem_ctrl_mem : wb_ctrl_mem;
  assign GEN_133 = T_7816 ? mem_ctrl_mem_cmd : wb_ctrl_mem_cmd;
  assign GEN_134 = T_7816 ? mem_ctrl_mem_type : wb_ctrl_mem_type;
  assign GEN_135 = T_7816 ? mem_ctrl_rfs1 : wb_ctrl_rfs1;
  assign GEN_136 = T_7816 ? mem_ctrl_rfs2 : wb_ctrl_rfs2;
  assign GEN_137 = T_7816 ? mem_ctrl_rfs3 : wb_ctrl_rfs3;
  assign GEN_138 = T_7816 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign GEN_139 = T_7816 ? mem_ctrl_div : wb_ctrl_div;
  assign GEN_140 = T_7816 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign GEN_141 = T_7816 ? mem_ctrl_csr : wb_ctrl_csr;
  assign GEN_142 = T_7816 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign GEN_143 = T_7816 ? mem_ctrl_fence : wb_ctrl_fence;
  assign GEN_144 = T_7816 ? mem_ctrl_amo : wb_ctrl_amo;
  assign GEN_145 = T_7816 ? T_7818 : wb_reg_wdata;
  assign GEN_146 = T_7816 ? GEN_118 : wb_reg_rs2;
  assign GEN_147 = T_7816 ? mem_reg_inst : wb_reg_inst;
  assign GEN_148 = T_7816 ? mem_reg_pc : wb_reg_pc;
  assign T_7819 = wb_ctrl_div | wb_dcache_miss;
  assign wb_set_sboard = T_7819 | wb_ctrl_rocc;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay;
  assign T_7822 = io_rocc_cmd_ready == 1'h0;
  assign T_7823 = T_7303 & T_7822;
  assign replay_wb = replay_wb_common | T_7823;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T_7824 = replay_wb | wb_xcpt;
  assign T_7825 = T_7824 | csr_io_eret;
  assign T_7826 = io_dmem_resp_bits_tag[0];
  assign dmem_resp_xpu = T_7826 == 1'h0;
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[8:1];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay;
  assign T_7830 = wb_reg_valid & wb_ctrl_wxd;
  assign T_7832 = T_7830 == 1'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign ll_waddr = GEN_150;
  assign T_7833 = div_io_resp_ready & div_io_resp_valid;
  assign ll_wen = GEN_151;
  assign T_7834 = dmem_resp_replay & dmem_resp_xpu;
  assign GEN_149 = T_7834 ? 1'h0 : T_7832;
  assign GEN_150 = T_7834 ? dmem_resp_waddr : {{3'd0}, div_io_resp_bits_tag};
  assign GEN_151 = T_7834 ? 1'h1 : T_7833;
  assign T_7838 = replay_wb == 1'h0;
  assign T_7839 = wb_reg_valid & T_7838;
  assign T_7841 = csr_io_csr_xcpt == 1'h0;
  assign wb_valid = T_7839 & T_7841;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign rf_wen = wb_wen | ll_wen;
  assign rf_waddr = ll_wen ? ll_waddr : {{3'd0}, wb_waddr};
  assign T_7842 = dmem_resp_valid & dmem_resp_xpu;
  assign T_7843 = wb_ctrl_csr != 3'h0;
  assign T_7844 = T_7843 ? csr_io_rw_rdata : wb_reg_wdata;
  assign T_7845 = ll_wen ? ll_wdata : T_7844;
  assign rf_wdata = T_7842 ? io_dmem_resp_bits_data : T_7845;
  assign GEN_195 = {{7'd0}, 1'h0};
  assign T_7847 = rf_waddr != GEN_195;
  assign T_7848 = rf_waddr[4:0];
  assign T_7849 = ~ T_7848;
  assign GEN_196 = {{3'd0}, id_raddr1};
  assign T_7851 = rf_waddr == GEN_196;
  assign GEN_152 = T_7851 ? rf_wdata : T_7194;
  assign GEN_197 = {{3'd0}, id_raddr2};
  assign T_7852 = rf_waddr == GEN_197;
  assign GEN_153 = T_7852 ? rf_wdata : T_7205;
  assign GEN_159 = T_7847 ? GEN_152 : T_7194;
  assign GEN_160 = T_7847 ? GEN_153 : T_7205;
  assign GEN_163 = rf_wen ? T_7847 : 1'h0;
  assign GEN_166 = rf_wen ? GEN_159 : T_7194;
  assign GEN_167 = rf_wen ? GEN_160 : T_7205;
  assign T_7853 = wb_reg_wdata[63:38];
  assign T_7854 = wb_reg_wdata[39:38];
  assign T_7855 = $signed(T_7854);
  assign T_7857 = T_7853 == GEN_183;
  assign T_7859 = T_7853 == GEN_184;
  assign T_7860 = T_7857 | T_7859;
  assign T_7862 = $signed(T_7855) != $signed(GEN_186);
  assign T_7863 = $signed(T_7853);
  assign T_7865 = $signed(T_7863) == $signed(GEN_188);
  assign T_7868 = $signed(T_7863) == $signed(GEN_190);
  assign T_7869 = T_7865 | T_7868;
  assign T_7871 = $signed(T_7855) == $signed(GEN_192);
  assign T_7872 = T_7855[0];
  assign T_7873 = T_7869 ? T_7871 : T_7872;
  assign T_7874 = T_7860 ? T_7862 : T_7873;
  assign T_7875 = wb_reg_wdata[38:0];
  assign T_7876 = {T_7874,T_7875};
  assign T_7877 = wb_reg_mem_xcpt ? T_7876 : wb_reg_pc;
  assign T_7894 = wb_reg_inst[31:20];
  assign T_7895 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T_7897 = id_raddr1 != GEN_170;
  assign T_7898 = id_ctrl_rxs1 & T_7897;
  assign T_7900 = id_raddr2 != GEN_170;
  assign T_7901 = id_ctrl_rxs2 & T_7900;
  assign T_7903 = id_waddr != GEN_170;
  assign T_7904 = id_ctrl_wxd & T_7903;
  assign GEN_211 = {{255'd0}, 1'h1};
  assign T_7909 = GEN_211 << ll_waddr;
  assign T_7911 = ll_wen ? T_7909 : {{255'd0}, 1'h0};
  assign T_7912 = ~ T_7911;
  assign GEN_212 = {{224'd0}, T_7906};
  assign T_7913 = GEN_212 & T_7912;
  assign GEN_168 = ll_wen ? T_7913 : {{224'd0}, T_7906};
  assign T_7915 = T_7906 >> id_raddr1;
  assign T_7916 = T_7915[0];
  assign T_7917 = T_7898 & T_7916;
  assign T_7918 = T_7906 >> id_raddr2;
  assign T_7919 = T_7918[0];
  assign T_7920 = T_7901 & T_7919;
  assign T_7921 = T_7906 >> id_waddr;
  assign T_7922 = T_7921[0];
  assign T_7923 = T_7904 & T_7922;
  assign T_7924 = T_7917 | T_7920;
  assign id_sboard_hazard = T_7924 | T_7923;
  assign T_7925 = wb_set_sboard & wb_wen;
  assign GEN_213 = {{31'd0}, 1'h1};
  assign T_7927 = GEN_213 << wb_waddr;
  assign T_7929 = T_7925 ? T_7927 : {{31'd0}, 1'h0};
  assign GEN_214 = {{224'd0}, T_7929};
  assign T_7930 = T_7913 | GEN_214;
  assign T_7931 = ll_wen | T_7925;
  assign GEN_169 = T_7931 ? T_7930 : GEN_168;
  assign T_7932 = ex_ctrl_csr != 3'h0;
  assign T_7933 = T_7932 | ex_ctrl_jalr;
  assign T_7934 = T_7933 | ex_ctrl_mem;
  assign T_7935 = T_7934 | ex_ctrl_div;
  assign T_7936 = T_7935 | ex_ctrl_fp;
  assign ex_cannot_bypass = T_7936 | ex_ctrl_rocc;
  assign T_7937 = id_raddr1 == ex_waddr;
  assign T_7938 = T_7898 & T_7937;
  assign T_7939 = id_raddr2 == ex_waddr;
  assign T_7940 = T_7901 & T_7939;
  assign T_7941 = id_waddr == ex_waddr;
  assign T_7942 = T_7904 & T_7941;
  assign T_7943 = T_7938 | T_7940;
  assign T_7944 = T_7943 | T_7942;
  assign data_hazard_ex = ex_ctrl_wxd & T_7944;
  assign T_7946 = io_fpu_dec_ren1 & T_7937;
  assign T_7948 = io_fpu_dec_ren2 & T_7939;
  assign T_7949 = id_raddr3 == ex_waddr;
  assign T_7950 = io_fpu_dec_ren3 & T_7949;
  assign T_7952 = io_fpu_dec_wen & T_7941;
  assign T_7953 = T_7946 | T_7948;
  assign T_7954 = T_7953 | T_7950;
  assign T_7955 = T_7954 | T_7952;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T_7955;
  assign T_7956 = data_hazard_ex & ex_cannot_bypass;
  assign T_7957 = T_7956 | fp_data_hazard_ex;
  assign id_ex_hazard = ex_reg_valid & T_7957;
  assign T_7959 = mem_ctrl_csr != 3'h0;
  assign T_7960 = mem_ctrl_mem & mem_reg_slow_bypass;
  assign T_7961 = T_7959 | T_7960;
  assign T_7962 = T_7961 | mem_ctrl_div;
  assign T_7963 = T_7962 | mem_ctrl_fp;
  assign mem_cannot_bypass = T_7963 | mem_ctrl_rocc;
  assign T_7964 = id_raddr1 == mem_waddr;
  assign T_7965 = T_7898 & T_7964;
  assign T_7966 = id_raddr2 == mem_waddr;
  assign T_7967 = T_7901 & T_7966;
  assign T_7968 = id_waddr == mem_waddr;
  assign T_7969 = T_7904 & T_7968;
  assign T_7970 = T_7965 | T_7967;
  assign T_7971 = T_7970 | T_7969;
  assign data_hazard_mem = mem_ctrl_wxd & T_7971;
  assign T_7973 = io_fpu_dec_ren1 & T_7964;
  assign T_7975 = io_fpu_dec_ren2 & T_7966;
  assign T_7976 = id_raddr3 == mem_waddr;
  assign T_7977 = io_fpu_dec_ren3 & T_7976;
  assign T_7979 = io_fpu_dec_wen & T_7968;
  assign T_7980 = T_7973 | T_7975;
  assign T_7981 = T_7980 | T_7977;
  assign T_7982 = T_7981 | T_7979;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T_7982;
  assign T_7983 = data_hazard_mem & mem_cannot_bypass;
  assign T_7984 = T_7983 | fp_data_hazard_mem;
  assign id_mem_hazard = mem_reg_valid & T_7984;
  assign T_7985 = mem_reg_valid & data_hazard_mem;
  assign T_7986 = T_7985 & mem_ctrl_mem;
  assign T_7987 = id_raddr1 == wb_waddr;
  assign T_7988 = T_7898 & T_7987;
  assign T_7989 = id_raddr2 == wb_waddr;
  assign T_7990 = T_7901 & T_7989;
  assign T_7991 = id_waddr == wb_waddr;
  assign T_7992 = T_7904 & T_7991;
  assign T_7993 = T_7988 | T_7990;
  assign T_7994 = T_7993 | T_7992;
  assign data_hazard_wb = wb_ctrl_wxd & T_7994;
  assign T_7996 = io_fpu_dec_ren1 & T_7987;
  assign T_7998 = io_fpu_dec_ren2 & T_7989;
  assign T_7999 = id_raddr3 == wb_waddr;
  assign T_8000 = io_fpu_dec_ren3 & T_7999;
  assign T_8002 = io_fpu_dec_wen & T_7991;
  assign T_8003 = T_7996 | T_7998;
  assign T_8004 = T_8003 | T_8000;
  assign T_8005 = T_8004 | T_8002;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T_8005;
  assign T_8006 = data_hazard_wb & wb_set_sboard;
  assign T_8007 = T_8006 | fp_data_hazard_wb;
  assign id_wb_hazard = wb_reg_valid & T_8007;
  assign T_8011 = io_dmem_req_valid | dcache_blocked;
  assign T_8012 = T_7516 & T_8011;
  assign T_8015 = wb_reg_xcpt == 1'h0;
  assign T_8018 = T_8015 & T_7822;
  assign T_8019 = io_rocc_cmd_valid | rocc_blocked;
  assign T_8020 = T_8018 & T_8019;
  assign T_8021 = id_ex_hazard | id_mem_hazard;
  assign T_8022 = T_8021 | id_wb_hazard;
  assign T_8023 = T_8022 | id_sboard_hazard;
  assign T_8026 = id_ctrl_mem & dcache_blocked;
  assign T_8027 = T_8023 | T_8026;
  assign T_8028 = id_ctrl_rocc & rocc_blocked;
  assign T_8029 = T_8027 | T_8028;
  assign T_8030 = T_8029 | T_7314;
  assign ctrl_stalld = T_8030 | csr_io_csr_stall;
  assign T_8032 = io_imem_resp_valid == 1'h0;
  assign T_8033 = T_8032 | take_pc_mem_wb;
  assign T_8034 = T_8033 | ctrl_stalld;
  assign T_8035 = T_8034 | csr_io_interrupt;
  assign T_8036 = wb_xcpt | csr_io_eret;
  assign T_8037 = replay_wb ? wb_reg_pc : mem_npc;
  assign T_8038 = T_8036 ? csr_io_evec : T_8037;
  assign T_8039 = wb_reg_valid & wb_ctrl_fence_i;
  assign T_8041 = io_dmem_s2_nack == 1'h0;
  assign T_8042 = T_8039 & T_8041;
  assign T_8044 = ctrl_stalld == 1'h0;
  assign T_8045 = T_8044 | csr_io_interrupt;
  assign T_8046 = T_8045 | take_pc_mem;
  assign T_8049 = mem_reg_valid & T_7732;
  assign T_8050 = T_8049 & mem_wrong_npc;
  assign T_8051 = T_8050 & mem_cfi_taken;
  assign T_8054 = T_8051 & T_7805;
  assign T_8055 = mem_ctrl_jal | mem_ctrl_jalr;
  assign T_8056 = mem_reg_inst[19:15];
  assign T_8059 = T_8056 & 5'h19;
  assign GEN_215 = {{4'd0}, 1'h1};
  assign T_8060 = GEN_215 == T_8059;
  assign T_8061 = mem_ctrl_jalr & T_8060;
  assign T_8062 = mem_reg_valid & mem_ctrl_branch;
  assign T_8065 = T_8062 & T_7805;
  assign T_8066 = mem_reg_valid & io_imem_btb_update_bits_isJump;
  assign T_8069 = T_8066 & T_7732;
  assign T_8072 = T_8069 & T_7805;
  assign T_8073 = mem_waddr[0];
  assign T_8074 = mem_ctrl_wxd & T_8073;
  assign T_8077 = T_7465 & id_ctrl_fp;
  assign T_8078 = dmem_resp_valid & T_7826;
  assign T_8079 = ex_reg_valid & ex_ctrl_mem;
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp};
  assign T_8081 = T_7375[63:38];
  assign T_8082 = alu_io_adder_out[39:38];
  assign T_8083 = $signed(T_8082);
  assign T_8085 = T_8081 == GEN_183;
  assign T_8087 = T_8081 == GEN_184;
  assign T_8088 = T_8085 | T_8087;
  assign T_8090 = $signed(T_8083) != $signed(GEN_186);
  assign T_8091 = $signed(T_8081);
  assign T_8093 = $signed(T_8091) == $signed(GEN_188);
  assign T_8096 = $signed(T_8091) == $signed(GEN_190);
  assign T_8097 = T_8093 | T_8096;
  assign T_8099 = $signed(T_8083) == $signed(GEN_192);
  assign T_8100 = T_8083[0];
  assign T_8101 = T_8097 ? T_8099 : T_8100;
  assign T_8102 = T_8088 ? T_8090 : T_8101;
  assign T_8103 = alu_io_adder_out[38:0];
  assign T_8104 = {T_8102,T_8103};
  assign T_8106 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign T_8109 = replay_wb_common == 1'h0;
  assign T_8110 = T_7303 & T_8109;
  assign T_8113 = wb_xcpt & T_7291;
  assign T_8132_funct = T_8150;
  assign T_8132_rs2 = T_8149;
  assign T_8132_rs1 = T_8148;
  assign T_8132_xd = T_8147;
  assign T_8132_xs1 = T_8146;
  assign T_8132_xs2 = T_8145;
  assign T_8132_rd = T_8144;
  assign T_8132_opcode = T_8143;
  assign T_8142 = wb_reg_inst;
  assign T_8143 = T_8142[6:0];
  assign T_8144 = T_8142[11:7];
  assign T_8145 = T_8142[12];
  assign T_8146 = T_8142[13];
  assign T_8147 = T_8142[14];
  assign T_8148 = T_8142[19:15];
  assign T_8149 = T_8142[24:20];
  assign T_8150 = T_8142[31:25];
  assign T_8151 = csr_io_time[31:0];
  assign T_8153 = rf_wen ? rf_waddr : {{7'd0}, 1'h0};
  assign T_8154 = wb_reg_inst[19:15];
  assign T_8157 = wb_reg_inst[24:20];
  assign T_8161 = reset == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_290 = {1{$random}};
  ex_ctrl_legal = GEN_290[0:0];
  GEN_291 = {1{$random}};
  ex_ctrl_fp = GEN_291[0:0];
  GEN_292 = {1{$random}};
  ex_ctrl_rocc = GEN_292[0:0];
  GEN_293 = {1{$random}};
  ex_ctrl_branch = GEN_293[0:0];
  GEN_294 = {1{$random}};
  ex_ctrl_jal = GEN_294[0:0];
  GEN_295 = {1{$random}};
  ex_ctrl_jalr = GEN_295[0:0];
  GEN_296 = {1{$random}};
  ex_ctrl_rxs2 = GEN_296[0:0];
  GEN_297 = {1{$random}};
  ex_ctrl_rxs1 = GEN_297[0:0];
  GEN_298 = {1{$random}};
  ex_ctrl_sel_alu2 = GEN_298[1:0];
  GEN_299 = {1{$random}};
  ex_ctrl_sel_alu1 = GEN_299[1:0];
  GEN_300 = {1{$random}};
  ex_ctrl_sel_imm = GEN_300[2:0];
  GEN_301 = {1{$random}};
  ex_ctrl_alu_dw = GEN_301[0:0];
  GEN_302 = {1{$random}};
  ex_ctrl_alu_fn = GEN_302[3:0];
  GEN_303 = {1{$random}};
  ex_ctrl_mem = GEN_303[0:0];
  GEN_304 = {1{$random}};
  ex_ctrl_mem_cmd = GEN_304[4:0];
  GEN_305 = {1{$random}};
  ex_ctrl_mem_type = GEN_305[2:0];
  GEN_306 = {1{$random}};
  ex_ctrl_rfs1 = GEN_306[0:0];
  GEN_307 = {1{$random}};
  ex_ctrl_rfs2 = GEN_307[0:0];
  GEN_308 = {1{$random}};
  ex_ctrl_rfs3 = GEN_308[0:0];
  GEN_309 = {1{$random}};
  ex_ctrl_wfd = GEN_309[0:0];
  GEN_310 = {1{$random}};
  ex_ctrl_div = GEN_310[0:0];
  GEN_311 = {1{$random}};
  ex_ctrl_wxd = GEN_311[0:0];
  GEN_312 = {1{$random}};
  ex_ctrl_csr = GEN_312[2:0];
  GEN_313 = {1{$random}};
  ex_ctrl_fence_i = GEN_313[0:0];
  GEN_314 = {1{$random}};
  ex_ctrl_fence = GEN_314[0:0];
  GEN_315 = {1{$random}};
  ex_ctrl_amo = GEN_315[0:0];
  GEN_316 = {1{$random}};
  mem_ctrl_legal = GEN_316[0:0];
  GEN_317 = {1{$random}};
  mem_ctrl_fp = GEN_317[0:0];
  GEN_318 = {1{$random}};
  mem_ctrl_rocc = GEN_318[0:0];
  GEN_319 = {1{$random}};
  mem_ctrl_branch = GEN_319[0:0];
  GEN_320 = {1{$random}};
  mem_ctrl_jal = GEN_320[0:0];
  GEN_321 = {1{$random}};
  mem_ctrl_jalr = GEN_321[0:0];
  GEN_322 = {1{$random}};
  mem_ctrl_rxs2 = GEN_322[0:0];
  GEN_323 = {1{$random}};
  mem_ctrl_rxs1 = GEN_323[0:0];
  GEN_324 = {1{$random}};
  mem_ctrl_sel_alu2 = GEN_324[1:0];
  GEN_325 = {1{$random}};
  mem_ctrl_sel_alu1 = GEN_325[1:0];
  GEN_326 = {1{$random}};
  mem_ctrl_sel_imm = GEN_326[2:0];
  GEN_327 = {1{$random}};
  mem_ctrl_alu_dw = GEN_327[0:0];
  GEN_328 = {1{$random}};
  mem_ctrl_alu_fn = GEN_328[3:0];
  GEN_329 = {1{$random}};
  mem_ctrl_mem = GEN_329[0:0];
  GEN_330 = {1{$random}};
  mem_ctrl_mem_cmd = GEN_330[4:0];
  GEN_331 = {1{$random}};
  mem_ctrl_mem_type = GEN_331[2:0];
  GEN_332 = {1{$random}};
  mem_ctrl_rfs1 = GEN_332[0:0];
  GEN_333 = {1{$random}};
  mem_ctrl_rfs2 = GEN_333[0:0];
  GEN_334 = {1{$random}};
  mem_ctrl_rfs3 = GEN_334[0:0];
  GEN_335 = {1{$random}};
  mem_ctrl_wfd = GEN_335[0:0];
  GEN_336 = {1{$random}};
  mem_ctrl_div = GEN_336[0:0];
  GEN_337 = {1{$random}};
  mem_ctrl_wxd = GEN_337[0:0];
  GEN_338 = {1{$random}};
  mem_ctrl_csr = GEN_338[2:0];
  GEN_339 = {1{$random}};
  mem_ctrl_fence_i = GEN_339[0:0];
  GEN_340 = {1{$random}};
  mem_ctrl_fence = GEN_340[0:0];
  GEN_341 = {1{$random}};
  mem_ctrl_amo = GEN_341[0:0];
  GEN_342 = {1{$random}};
  wb_ctrl_legal = GEN_342[0:0];
  GEN_343 = {1{$random}};
  wb_ctrl_fp = GEN_343[0:0];
  GEN_344 = {1{$random}};
  wb_ctrl_rocc = GEN_344[0:0];
  GEN_345 = {1{$random}};
  wb_ctrl_branch = GEN_345[0:0];
  GEN_346 = {1{$random}};
  wb_ctrl_jal = GEN_346[0:0];
  GEN_347 = {1{$random}};
  wb_ctrl_jalr = GEN_347[0:0];
  GEN_348 = {1{$random}};
  wb_ctrl_rxs2 = GEN_348[0:0];
  GEN_349 = {1{$random}};
  wb_ctrl_rxs1 = GEN_349[0:0];
  GEN_350 = {1{$random}};
  wb_ctrl_sel_alu2 = GEN_350[1:0];
  GEN_351 = {1{$random}};
  wb_ctrl_sel_alu1 = GEN_351[1:0];
  GEN_352 = {1{$random}};
  wb_ctrl_sel_imm = GEN_352[2:0];
  GEN_353 = {1{$random}};
  wb_ctrl_alu_dw = GEN_353[0:0];
  GEN_354 = {1{$random}};
  wb_ctrl_alu_fn = GEN_354[3:0];
  GEN_355 = {1{$random}};
  wb_ctrl_mem = GEN_355[0:0];
  GEN_356 = {1{$random}};
  wb_ctrl_mem_cmd = GEN_356[4:0];
  GEN_357 = {1{$random}};
  wb_ctrl_mem_type = GEN_357[2:0];
  GEN_358 = {1{$random}};
  wb_ctrl_rfs1 = GEN_358[0:0];
  GEN_359 = {1{$random}};
  wb_ctrl_rfs2 = GEN_359[0:0];
  GEN_360 = {1{$random}};
  wb_ctrl_rfs3 = GEN_360[0:0];
  GEN_361 = {1{$random}};
  wb_ctrl_wfd = GEN_361[0:0];
  GEN_362 = {1{$random}};
  wb_ctrl_div = GEN_362[0:0];
  GEN_363 = {1{$random}};
  wb_ctrl_wxd = GEN_363[0:0];
  GEN_364 = {1{$random}};
  wb_ctrl_csr = GEN_364[2:0];
  GEN_365 = {1{$random}};
  wb_ctrl_fence_i = GEN_365[0:0];
  GEN_366 = {1{$random}};
  wb_ctrl_fence = GEN_366[0:0];
  GEN_367 = {1{$random}};
  wb_ctrl_amo = GEN_367[0:0];
  GEN_368 = {1{$random}};
  ex_reg_xcpt_interrupt = GEN_368[0:0];
  GEN_369 = {1{$random}};
  ex_reg_valid = GEN_369[0:0];
  GEN_370 = {1{$random}};
  ex_reg_btb_hit = GEN_370[0:0];
  GEN_371 = {1{$random}};
  ex_reg_btb_resp_taken = GEN_371[0:0];
  GEN_372 = {1{$random}};
  ex_reg_btb_resp_mask = GEN_372[0:0];
  GEN_373 = {1{$random}};
  ex_reg_btb_resp_bridx = GEN_373[0:0];
  GEN_374 = {2{$random}};
  ex_reg_btb_resp_target = GEN_374[38:0];
  GEN_375 = {1{$random}};
  ex_reg_btb_resp_entry = GEN_375[5:0];
  GEN_376 = {1{$random}};
  ex_reg_btb_resp_bht_history = GEN_376[6:0];
  GEN_377 = {1{$random}};
  ex_reg_btb_resp_bht_value = GEN_377[1:0];
  GEN_378 = {1{$random}};
  ex_reg_xcpt = GEN_378[0:0];
  GEN_379 = {1{$random}};
  ex_reg_flush_pipe = GEN_379[0:0];
  GEN_380 = {1{$random}};
  ex_reg_load_use = GEN_380[0:0];
  GEN_381 = {2{$random}};
  ex_reg_cause = GEN_381[63:0];
  GEN_382 = {2{$random}};
  ex_reg_pc = GEN_382[39:0];
  GEN_383 = {1{$random}};
  ex_reg_inst = GEN_383[31:0];
  GEN_384 = {1{$random}};
  mem_reg_xcpt_interrupt = GEN_384[0:0];
  GEN_385 = {1{$random}};
  mem_reg_valid = GEN_385[0:0];
  GEN_386 = {1{$random}};
  mem_reg_btb_hit = GEN_386[0:0];
  GEN_387 = {1{$random}};
  mem_reg_btb_resp_taken = GEN_387[0:0];
  GEN_388 = {1{$random}};
  mem_reg_btb_resp_mask = GEN_388[0:0];
  GEN_389 = {1{$random}};
  mem_reg_btb_resp_bridx = GEN_389[0:0];
  GEN_390 = {2{$random}};
  mem_reg_btb_resp_target = GEN_390[38:0];
  GEN_391 = {1{$random}};
  mem_reg_btb_resp_entry = GEN_391[5:0];
  GEN_392 = {1{$random}};
  mem_reg_btb_resp_bht_history = GEN_392[6:0];
  GEN_393 = {1{$random}};
  mem_reg_btb_resp_bht_value = GEN_393[1:0];
  GEN_394 = {1{$random}};
  mem_reg_xcpt = GEN_394[0:0];
  GEN_395 = {1{$random}};
  mem_reg_replay = GEN_395[0:0];
  GEN_396 = {1{$random}};
  mem_reg_flush_pipe = GEN_396[0:0];
  GEN_397 = {2{$random}};
  mem_reg_cause = GEN_397[63:0];
  GEN_398 = {1{$random}};
  mem_reg_slow_bypass = GEN_398[0:0];
  GEN_399 = {1{$random}};
  mem_reg_load = GEN_399[0:0];
  GEN_400 = {1{$random}};
  mem_reg_store = GEN_400[0:0];
  GEN_401 = {2{$random}};
  mem_reg_pc = GEN_401[39:0];
  GEN_402 = {1{$random}};
  mem_reg_inst = GEN_402[31:0];
  GEN_403 = {2{$random}};
  mem_reg_wdata = GEN_403[63:0];
  GEN_404 = {2{$random}};
  mem_reg_rs2 = GEN_404[63:0];
  GEN_405 = {1{$random}};
  wb_reg_valid = GEN_405[0:0];
  GEN_406 = {1{$random}};
  wb_reg_xcpt = GEN_406[0:0];
  GEN_407 = {1{$random}};
  wb_reg_mem_xcpt = GEN_407[0:0];
  GEN_408 = {1{$random}};
  wb_reg_replay = GEN_408[0:0];
  GEN_409 = {2{$random}};
  wb_reg_cause = GEN_409[63:0];
  GEN_410 = {2{$random}};
  wb_reg_pc = GEN_410[39:0];
  GEN_411 = {1{$random}};
  wb_reg_inst = GEN_411[31:0];
  GEN_412 = {2{$random}};
  wb_reg_wdata = GEN_412[63:0];
  GEN_413 = {2{$random}};
  wb_reg_rs2 = GEN_413[63:0];
  GEN_414 = {1{$random}};
  id_reg_fence = GEN_414[0:0];
  GEN_415 = {2{$random}};
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    T_7183[initvar] = GEN_415[63:0];
  GEN_416 = {1{$random}};
  ex_reg_rs_bypass_0 = GEN_416[0:0];
  GEN_417 = {1{$random}};
  ex_reg_rs_bypass_1 = GEN_417[0:0];
  GEN_418 = {1{$random}};
  ex_reg_rs_lsb_0 = GEN_418[1:0];
  GEN_419 = {1{$random}};
  ex_reg_rs_lsb_1 = GEN_419[1:0];
  GEN_420 = {2{$random}};
  ex_reg_rs_msb_0 = GEN_420[61:0];
  GEN_421 = {2{$random}};
  ex_reg_rs_msb_1 = GEN_421[61:0];
  GEN_422 = {1{$random}};
  T_7799 = GEN_422[0:0];
  GEN_423 = {1{$random}};
  T_7906 = GEN_423[31:0];
  GEN_424 = {1{$random}};
  dcache_blocked = GEN_424[0:0];
  GEN_425 = {1{$random}};
  rocc_blocked = GEN_425[0:0];
  GEN_426 = {2{$random}};
  T_8155 = GEN_426[63:0];
  GEN_427 = {2{$random}};
  T_8156 = GEN_427[63:0];
  GEN_428 = {2{$random}};
  T_8158 = GEN_428[63:0];
  GEN_429 = {2{$random}};
  T_8159 = GEN_429[63:0];
  GEN_430 = {1{$random}};
  GEN_154 = GEN_430[0:0];
  GEN_431 = {2{$random}};
  GEN_155 = GEN_431[63:0];
  GEN_432 = {1{$random}};
  GEN_156 = GEN_432[0:0];
  GEN_433 = {1{$random}};
  GEN_157 = GEN_433[4:0];
  GEN_434 = {1{$random}};
  GEN_158 = GEN_434[0:0];
  GEN_435 = {1{$random}};
  GEN_161 = GEN_435[0:0];
  GEN_436 = {1{$random}};
  GEN_162 = GEN_436[0:0];
  GEN_437 = {1{$random}};
  GEN_164 = GEN_437[0:0];
  GEN_438 = {1{$random}};
  GEN_165 = GEN_438[0:0];
  GEN_439 = {1{$random}};
  GEN_171 = GEN_439[0:0];
  GEN_440 = {1{$random}};
  GEN_172 = GEN_440[0:0];
  GEN_441 = {1{$random}};
  GEN_174 = GEN_441[0:0];
  GEN_442 = {1{$random}};
  GEN_175 = GEN_442[0:0];
  GEN_443 = {1{$random}};
  GEN_176 = GEN_443[0:0];
  GEN_444 = {1{$random}};
  GEN_178 = GEN_444[0:0];
  GEN_445 = {1{$random}};
  GEN_180 = GEN_445[0:0];
  GEN_446 = {1{$random}};
  GEN_185 = GEN_446[0:0];
  GEN_447 = {1{$random}};
  GEN_191 = GEN_447[0:0];
  GEN_448 = {1{$random}};
  GEN_193 = GEN_448[0:0];
  GEN_449 = {1{$random}};
  GEN_198 = GEN_449[0:0];
  GEN_450 = {1{$random}};
  GEN_199 = GEN_450[2:0];
  GEN_451 = {1{$random}};
  GEN_200 = GEN_451[1:0];
  GEN_452 = {3{$random}};
  GEN_201 = GEN_452[64:0];
  GEN_453 = {3{$random}};
  GEN_202 = GEN_453[64:0];
  GEN_454 = {3{$random}};
  GEN_203 = GEN_454[64:0];
  GEN_455 = {1{$random}};
  GEN_204 = GEN_455[0:0];
  GEN_456 = {1{$random}};
  GEN_205 = GEN_456[0:0];
  GEN_457 = {1{$random}};
  GEN_206 = GEN_457[0:0];
  GEN_458 = {1{$random}};
  GEN_207 = GEN_458[0:0];
  GEN_459 = {1{$random}};
  GEN_208 = GEN_459[0:0];
  GEN_460 = {2{$random}};
  GEN_209 = GEN_460[39:0];
  GEN_461 = {1{$random}};
  GEN_210 = GEN_461[8:0];
  GEN_462 = {1{$random}};
  GEN_216 = GEN_462[4:0];
  GEN_463 = {1{$random}};
  GEN_217 = GEN_463[2:0];
  GEN_464 = {2{$random}};
  GEN_218 = GEN_464[63:0];
  GEN_465 = {1{$random}};
  GEN_219 = GEN_465[0:0];
  GEN_466 = {1{$random}};
  GEN_220 = GEN_466[0:0];
  GEN_467 = {2{$random}};
  GEN_221 = GEN_467[63:0];
  GEN_468 = {2{$random}};
  GEN_222 = GEN_468[63:0];
  GEN_469 = {1{$random}};
  GEN_223 = GEN_469[0:0];
  GEN_470 = {1{$random}};
  GEN_224 = GEN_470[0:0];
  GEN_471 = {1{$random}};
  GEN_225 = GEN_471[0:0];
  GEN_472 = {1{$random}};
  GEN_226 = GEN_472[0:0];
  GEN_473 = {1{$random}};
  GEN_227 = GEN_473[0:0];
  GEN_474 = {1{$random}};
  GEN_228 = GEN_474[0:0];
  GEN_475 = {1{$random}};
  GEN_229 = GEN_475[0:0];
  GEN_476 = {1{$random}};
  GEN_230 = GEN_476[0:0];
  GEN_477 = {1{$random}};
  GEN_231 = GEN_477[2:0];
  GEN_478 = {1{$random}};
  GEN_232 = GEN_478[1:0];
  GEN_479 = {1{$random}};
  GEN_233 = GEN_479[2:0];
  GEN_480 = {1{$random}};
  GEN_234 = GEN_480[0:0];
  GEN_481 = {1{$random}};
  GEN_235 = GEN_481[3:0];
  GEN_482 = {2{$random}};
  GEN_236 = GEN_482[63:0];
  GEN_483 = {1{$random}};
  GEN_237 = GEN_483[0:0];
  GEN_484 = {1{$random}};
  GEN_238 = GEN_484[0:0];
  GEN_485 = {3{$random}};
  GEN_239 = GEN_485[64:0];
  GEN_486 = {1{$random}};
  GEN_240 = GEN_486[4:0];
  GEN_487 = {1{$random}};
  GEN_241 = GEN_487[0:0];
  GEN_488 = {1{$random}};
  GEN_242 = GEN_488[0:0];
  GEN_489 = {1{$random}};
  GEN_243 = GEN_489[0:0];
  GEN_490 = {1{$random}};
  GEN_244 = GEN_490[4:0];
  GEN_491 = {2{$random}};
  GEN_245 = GEN_491[63:0];
  GEN_492 = {1{$random}};
  GEN_246 = GEN_492[0:0];
  GEN_493 = {2{$random}};
  GEN_247 = GEN_493[39:0];
  GEN_494 = {1{$random}};
  GEN_248 = GEN_494[8:0];
  GEN_495 = {1{$random}};
  GEN_249 = GEN_495[4:0];
  GEN_496 = {1{$random}};
  GEN_250 = GEN_496[2:0];
  GEN_497 = {1{$random}};
  GEN_251 = GEN_497[0:0];
  GEN_498 = {2{$random}};
  GEN_252 = GEN_498[63:0];
  GEN_499 = {1{$random}};
  GEN_253 = GEN_499[0:0];
  GEN_500 = {2{$random}};
  GEN_254 = GEN_500[63:0];
  GEN_501 = {1{$random}};
  GEN_255 = GEN_501[0:0];
  GEN_502 = {1{$random}};
  GEN_256 = GEN_502[0:0];
  GEN_503 = {1{$random}};
  GEN_257 = GEN_503[0:0];
  GEN_504 = {1{$random}};
  GEN_258 = GEN_504[25:0];
  GEN_505 = {1{$random}};
  GEN_259 = GEN_505[1:0];
  GEN_506 = {1{$random}};
  GEN_260 = GEN_506[2:0];
  GEN_507 = {1{$random}};
  GEN_261 = GEN_507[0:0];
  GEN_508 = {1{$random}};
  GEN_262 = GEN_508[2:0];
  GEN_509 = {1{$random}};
  GEN_263 = GEN_509[11:0];
  GEN_510 = {2{$random}};
  GEN_264 = GEN_510[63:0];
  GEN_511 = {1{$random}};
  GEN_265 = GEN_511[0:0];
  GEN_512 = {1{$random}};
  GEN_266 = GEN_512[0:0];
  GEN_513 = {1{$random}};
  GEN_267 = GEN_513[4:0];
  GEN_514 = {1{$random}};
  GEN_268 = GEN_514[0:0];
  GEN_515 = {1{$random}};
  GEN_269 = GEN_515[0:0];
  GEN_516 = {1{$random}};
  GEN_270 = GEN_516[0:0];
  GEN_517 = {1{$random}};
  GEN_271 = GEN_517[0:0];
  GEN_518 = {1{$random}};
  GEN_272 = GEN_518[0:0];
  GEN_519 = {1{$random}};
  GEN_273 = GEN_519[0:0];
  GEN_520 = {1{$random}};
  GEN_274 = GEN_520[0:0];
  GEN_521 = {1{$random}};
  GEN_275 = GEN_521[0:0];
  GEN_522 = {1{$random}};
  GEN_276 = GEN_522[0:0];
  GEN_523 = {1{$random}};
  GEN_277 = GEN_523[0:0];
  GEN_524 = {1{$random}};
  GEN_278 = GEN_524[0:0];
  GEN_525 = {1{$random}};
  GEN_279 = GEN_525[0:0];
  GEN_526 = {1{$random}};
  GEN_280 = GEN_526[0:0];
  GEN_527 = {1{$random}};
  GEN_281 = GEN_527[0:0];
  GEN_528 = {1{$random}};
  GEN_282 = GEN_528[0:0];
  GEN_529 = {1{$random}};
  GEN_283 = GEN_529[0:0];
  GEN_530 = {1{$random}};
  GEN_284 = GEN_530[2:0];
  GEN_531 = {1{$random}};
  GEN_285 = GEN_531[1:0];
  GEN_532 = {3{$random}};
  GEN_286 = GEN_532[64:0];
  GEN_533 = {3{$random}};
  GEN_287 = GEN_533[64:0];
  GEN_534 = {3{$random}};
  GEN_288 = GEN_534[64:0];
  GEN_535 = {1{$random}};
  GEN_289 = GEN_535[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_legal <= id_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_fp <= id_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_rocc <= id_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_branch <= id_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_jal <= id_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_jalr <= id_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_rxs2 <= id_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_rxs1 <= id_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_sel_imm <= id_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_alu_dw <= id_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_alu_fn <= id_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_mem <= id_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_mem_type <= id_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_rfs1 <= id_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_rfs2 <= id_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_rfs3 <= id_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_wfd <= id_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_div <= id_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_wxd <= id_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(id_csr_ren) begin
          ex_ctrl_csr <= 3'h5;
        end else begin
          ex_ctrl_csr <= id_ctrl_csr;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(T_7477) begin
          ex_ctrl_fence_i <= 1'h1;
        end else begin
          ex_ctrl_fence_i <= id_ctrl_fence_i;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_fence <= id_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_ctrl_amo <= id_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_legal <= ex_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fp <= ex_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rocc <= ex_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_branch <= ex_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_jal <= ex_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_jalr <= ex_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rxs2 <= ex_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rxs1 <= ex_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_alu2 <= ex_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_alu1 <= ex_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_imm <= ex_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_alu_dw <= ex_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_alu_fn <= ex_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem <= ex_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem_cmd <= ex_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem_type <= ex_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs1 <= ex_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs2 <= ex_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs3 <= ex_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_wfd <= ex_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_div <= ex_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_wxd <= ex_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_csr <= ex_ctrl_csr;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fence_i <= ex_ctrl_fence_i;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fence <= ex_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_amo <= ex_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_legal <= mem_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_fp <= mem_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_rocc <= mem_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_branch <= mem_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_jal <= mem_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_jalr <= mem_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_rxs2 <= mem_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_rxs1 <= mem_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_sel_alu2 <= mem_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_sel_alu1 <= mem_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_sel_imm <= mem_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_alu_dw <= mem_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_alu_fn <= mem_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_mem <= mem_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_mem_cmd <= mem_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_mem_type <= mem_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_rfs1 <= mem_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_rfs2 <= mem_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_rfs3 <= mem_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_wfd <= mem_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_div <= mem_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_wxd <= mem_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_csr <= mem_ctrl_csr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_fence_i <= mem_ctrl_fence_i;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_fence <= mem_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_ctrl_amo <= mem_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt_interrupt <= T_7472;
    end
    if(1'h0) begin
    end else begin
      ex_reg_valid <= T_7465;
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_reg_btb_hit <= io_imem_btb_resp_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_mask <= io_imem_btb_resp_bits_mask;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_bridx <= io_imem_btb_resp_bits_bridx;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
        end
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt <= T_7468;
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(T_7477) begin
          ex_reg_flush_pipe <= 1'h1;
        end else begin
          ex_reg_flush_pipe <= T_7476;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_reg_load_use <= id_load_use;
      end
    end
    if(1'h0) begin
    end else begin
      if(id_xcpt) begin
        if(csr_io_interrupt) begin
          ex_reg_cause <= csr_io_interrupt_cause;
        end else begin
          ex_reg_cause <= {{62'd0}, T_7321};
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7512) begin
        ex_reg_pc <= io_imem_resp_bits_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7512) begin
        ex_reg_inst <= io_imem_resp_bits_data_0;
      end
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt_interrupt <= T_7744;
    end
    if(1'h0) begin
    end else begin
      mem_reg_valid <= T_7735;
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_btb_hit <= ex_reg_btb_hit;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
        end
      end
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt <= T_7741;
    end
    if(1'h0) begin
    end else begin
      mem_reg_replay <= T_7738;
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_flush_pipe <= ex_reg_flush_pipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_xcpt) begin
        if(T_7542) begin
          mem_reg_cause <= ex_reg_cause;
        end else begin
          mem_reg_cause <= {{62'd0}, 2'h2};
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_slow_bypass <= ex_slow_bypass;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_load <= T_7754;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_store <= T_7762;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_pc <= ex_reg_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_wdata <= alu_io_out;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(T_7764) begin
          if(ex_reg_rs_bypass_1) begin
            mem_reg_rs2 <= GEN_1;
          end else begin
            mem_reg_rs2 <= T_7376;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      wb_reg_valid <= T_7803;
    end
    if(1'h0) begin
    end else begin
      wb_reg_xcpt <= T_7809;
    end
    if(1'h0) begin
    end else begin
      wb_reg_mem_xcpt <= T_7814;
    end
    if(1'h0) begin
    end else begin
      wb_reg_replay <= T_7806;
    end
    if(1'h0) begin
    end else begin
      if(mem_xcpt) begin
        if(T_7789) begin
          wb_reg_cause <= mem_reg_cause;
        end else begin
          wb_reg_cause <= {{61'd0}, mem_new_cause};
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_reg_pc <= mem_reg_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        wb_reg_inst <= mem_reg_inst;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        if(T_7817) begin
          wb_reg_wdata <= io_fpu_toint_data;
        end else begin
          wb_reg_wdata <= mem_int_wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7816) begin
        if(mem_ctrl_rocc) begin
          wb_reg_rs2 <= mem_reg_rs2;
        end
      end
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T_7306;
    end
    if(T_7183_T_7850_en & T_7183_T_7850_mask) begin
      T_7183[T_7183_T_7850_addr] <= T_7183_T_7850_data;
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_reg_rs_bypass_0 <= T_7482;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        ex_reg_rs_bypass_1 <= T_7497;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(T_7492) begin
          ex_reg_rs_lsb_0 <= T_7493;
        end else begin
          if(T_7331) begin
            ex_reg_rs_lsb_0 <= {{1'd0}, 1'h0};
          end else begin
            if(T_7334) begin
              ex_reg_rs_lsb_0 <= {{1'd0}, 1'h1};
            end else begin
              if(T_7336) begin
                ex_reg_rs_lsb_0 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_0 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(T_7507) begin
          ex_reg_rs_lsb_1 <= T_7508;
        end else begin
          if(T_7339) begin
            ex_reg_rs_lsb_1 <= {{1'd0}, 1'h0};
          end else begin
            if(T_7342) begin
              ex_reg_rs_lsb_1 <= {{1'd0}, 1'h1};
            end else begin
              if(T_7344) begin
                ex_reg_rs_lsb_1 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_1 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(T_7492) begin
          ex_reg_rs_msb_0 <= T_7494;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7465) begin
        if(T_7507) begin
          ex_reg_rs_msb_1 <= T_7509;
        end
      end
    end
    if(1'h0) begin
    end else begin
      T_7799 <= T_7798;
    end
    if(reset) begin
      T_7906 <= 32'h0;
    end else begin
      T_7906 <= GEN_169[31:0];
    end
    if(1'h0) begin
    end else begin
      dcache_blocked <= T_8012;
    end
    if(1'h0) begin
    end else begin
      rocc_blocked <= T_8020;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_rs_bypass_0) begin
        T_8155 <= GEN_0;
      end else begin
        T_8155 <= T_7374;
      end
    end
    if(1'h0) begin
    end else begin
      T_8156 <= T_8155;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_rs_bypass_1) begin
        T_8158 <= GEN_1;
      end else begin
        T_8158 <= T_7376;
      end
    end
    if(1'h0) begin
    end else begin
      T_8159 <= T_8158;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_8161) begin
          $fwrite(32'h80000002,"C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n",io_prci_id,T_8151,wb_valid,wb_reg_pc,T_8153,rf_wdata,rf_wen,T_8154,T_8156,T_8157,T_8159,wb_reg_inst,wb_reg_inst);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module FlowThroughSerializer(
  input   clk,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input  [2:0] io_in_bits_addr_beat,
  input  [1:0] io_in_bits_client_xact_id,
  input  [2:0] io_in_bits_manager_xact_id,
  input   io_in_bits_is_builtin_type,
  input  [3:0] io_in_bits_g_type,
  input  [63:0] io_in_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_cnt,
  output  io_done
);
  assign io_in_ready = io_out_ready;
  assign io_out_valid = io_in_valid;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_data = io_in_bits_data;
  assign io_cnt = 1'h0;
  assign io_done = 1'h1;
endmodule
module ICache(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [38:0] io_req_bits_addr,
  input  [19:0] io_s1_ppn,
  input   io_s1_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [31:0] io_resp_bits_data,
  output [63:0] io_resp_bits_datablock,
  input   io_invalidate,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  reg [1:0] state;
  reg [31:0] GEN_5;
  reg  invalidated;
  reg [31:0] GEN_6;
  wire  stall;
  wire  rdy;
  reg [31:0] refill_addr;
  reg [31:0] GEN_7;
  wire  s1_any_tag_hit;
  reg  s1_valid;
  reg [31:0] GEN_8;
  reg [38:0] s1_vaddr;
  reg [63:0] GEN_9;
  wire [11:0] T_934;
  wire [31:0] s1_paddr;
  wire [19:0] s1_tag;
  wire  T_935;
  wire [38:0] s0_vaddr;
  wire  T_937;
  wire  T_940;
  wire  T_941;
  wire  T_942;
  wire [38:0] GEN_0;
  wire  T_946;
  wire  T_947;
  wire  out_valid;
  wire [5:0] s1_idx;
  wire  s1_hit;
  wire  T_949;
  wire  s1_miss;
  wire  T_952;
  wire  T_953;
  wire  T_955;
  wire  T_956;
  wire [31:0] GEN_1;
  wire [19:0] refill_tag;
  wire  FlowThroughSerializer_1_clk;
  wire  FlowThroughSerializer_1_reset;
  wire  FlowThroughSerializer_1_io_in_ready;
  wire  FlowThroughSerializer_1_io_in_valid;
  wire [2:0] FlowThroughSerializer_1_io_in_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_1_io_in_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_1_io_in_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_io_in_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_io_in_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_io_in_bits_data;
  wire  FlowThroughSerializer_1_io_out_ready;
  wire  FlowThroughSerializer_1_io_out_valid;
  wire [2:0] FlowThroughSerializer_1_io_out_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_1_io_out_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_1_io_out_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_io_out_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_io_out_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_io_out_bits_data;
  wire  FlowThroughSerializer_1_io_cnt;
  wire  FlowThroughSerializer_1_io_done;
  wire  T_957;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_10;
  wire  T_960;
  wire [2:0] GEN_72;
  wire [3:0] T_962;
  wire [2:0] T_963;
  wire [2:0] GEN_2;
  wire  refill_wrap;
  wire  T_964;
  wire  refill_done;
  reg [15:0] T_967;
  reg [31:0] GEN_11;
  wire  T_968;
  wire  T_969;
  wire  T_970;
  wire  T_971;
  wire  T_972;
  wire  T_973;
  wire  T_974;
  wire [14:0] T_975;
  wire [15:0] T_976;
  wire [15:0] GEN_3;
  wire [1:0] repl_way;
  reg [19:0] tag_array_0 [0:63];
  reg [31:0] GEN_12;
  wire [19:0] tag_array_0_tag_rdata_data;
  wire [5:0] tag_array_0_tag_rdata_addr;
  wire  tag_array_0_tag_rdata_en;
  reg [5:0] GEN_13;
  reg [31:0] GEN_14;
  reg  GEN_15;
  reg [31:0] GEN_16;
  wire [19:0] tag_array_0_T_1018_data;
  wire [5:0] tag_array_0_T_1018_addr;
  wire  tag_array_0_T_1018_mask;
  wire  tag_array_0_T_1018_en;
  reg [19:0] tag_array_1 [0:63];
  reg [31:0] GEN_17;
  wire [19:0] tag_array_1_tag_rdata_data;
  wire [5:0] tag_array_1_tag_rdata_addr;
  wire  tag_array_1_tag_rdata_en;
  reg [5:0] GEN_18;
  reg [31:0] GEN_19;
  reg  GEN_20;
  reg [31:0] GEN_21;
  wire [19:0] tag_array_1_T_1018_data;
  wire [5:0] tag_array_1_T_1018_addr;
  wire  tag_array_1_T_1018_mask;
  wire  tag_array_1_T_1018_en;
  reg [19:0] tag_array_2 [0:63];
  reg [31:0] GEN_22;
  wire [19:0] tag_array_2_tag_rdata_data;
  wire [5:0] tag_array_2_tag_rdata_addr;
  wire  tag_array_2_tag_rdata_en;
  reg [5:0] GEN_23;
  reg [31:0] GEN_24;
  reg  GEN_26;
  reg [31:0] GEN_28;
  wire [19:0] tag_array_2_T_1018_data;
  wire [5:0] tag_array_2_T_1018_addr;
  wire  tag_array_2_T_1018_mask;
  wire  tag_array_2_T_1018_en;
  reg [19:0] tag_array_3 [0:63];
  reg [31:0] GEN_30;
  wire [19:0] tag_array_3_tag_rdata_data;
  wire [5:0] tag_array_3_tag_rdata_addr;
  wire  tag_array_3_tag_rdata_en;
  reg [5:0] GEN_39;
  reg [31:0] GEN_40;
  reg  GEN_41;
  reg [31:0] GEN_43;
  wire [19:0] tag_array_3_T_1018_data;
  wire [5:0] tag_array_3_T_1018_addr;
  wire  tag_array_3_T_1018_mask;
  wire  tag_array_3_T_1018_en;
  wire [5:0] T_985;
  wire [5:0] T_990;
  wire [19:0] T_999_0;
  wire [19:0] T_999_1;
  wire [19:0] T_999_2;
  wire [19:0] T_999_3;
  wire [1:0] GEN_73;
  wire  T_1002;
  wire [1:0] GEN_74;
  wire  T_1004;
  wire  T_1006;
  wire  T_1008;
  wire  T_1014_0;
  wire  T_1014_1;
  wire  T_1014_2;
  wire  T_1014_3;
  wire  GEN_25;
  wire  GEN_27;
  wire  GEN_29;
  wire  GEN_31;
  reg [255:0] vb_array;
  reg [255:0] GEN_44;
  wire  T_1022;
  wire  T_1023;
  wire [7:0] T_1024;
  wire [255:0] GEN_75;
  wire [255:0] T_1027;
  wire [255:0] T_1028;
  wire [255:0] T_1029;
  wire [255:0] GEN_32;
  wire [255:0] GEN_33;
  wire  GEN_34;
  wire  s1_disparity_0;
  wire  s1_disparity_1;
  wire  s1_disparity_2;
  wire  s1_disparity_3;
  wire  T_1042;
  wire [6:0] T_1044;
  wire [127:0] GEN_76;
  wire [127:0] T_1047;
  wire [255:0] GEN_77;
  wire [255:0] T_1050;
  wire [255:0] T_1051;
  wire [255:0] GEN_35;
  wire  T_1053;
  wire [6:0] T_1055;
  wire [127:0] T_1058;
  wire [255:0] GEN_80;
  wire [255:0] T_1061;
  wire [255:0] T_1062;
  wire [255:0] GEN_36;
  wire  T_1064;
  wire [7:0] T_1066;
  wire [255:0] T_1069;
  wire [255:0] T_1072;
  wire [255:0] T_1073;
  wire [255:0] GEN_37;
  wire  T_1075;
  wire [7:0] T_1077;
  wire [255:0] T_1080;
  wire [255:0] T_1083;
  wire [255:0] T_1084;
  wire [255:0] GEN_38;
  wire  s1_tag_match_0;
  wire  s1_tag_match_1;
  wire  s1_tag_match_2;
  wire  s1_tag_match_3;
  wire  s1_tag_hit_0;
  wire  s1_tag_hit_1;
  wire  s1_tag_hit_2;
  wire  s1_tag_hit_3;
  wire [63:0] s1_dout_0;
  wire [63:0] s1_dout_1;
  wire [63:0] s1_dout_2;
  wire [63:0] s1_dout_3;
  wire  T_1108;
  wire [255:0] T_1112;
  wire  T_1113;
  wire  T_1115;
  wire [19:0] T_1119;
  wire  T_1120;
  wire  T_1121;
  wire [255:0] T_1132;
  wire  T_1133;
  wire  T_1135;
  wire [19:0] T_1139;
  wire  T_1140;
  wire  T_1141;
  wire [255:0] T_1152;
  wire  T_1153;
  wire  T_1155;
  wire [19:0] T_1159;
  wire  T_1160;
  wire  T_1161;
  wire [255:0] T_1172;
  wire  T_1173;
  wire  T_1175;
  wire [19:0] T_1179;
  wire  T_1180;
  wire  T_1181;
  wire  T_1187;
  wire  T_1188;
  wire  T_1189;
  wire  T_1190;
  wire  T_1191;
  wire  T_1192;
  wire  T_1194;
  wire  T_1195;
  reg [63:0] T_1198 [0:511];
  reg [63:0] GEN_45;
  wire [63:0] T_1198_T_1210_data;
  wire [8:0] T_1198_T_1210_addr;
  wire  T_1198_T_1210_en;
  reg [8:0] GEN_46;
  reg [31:0] GEN_47;
  reg  GEN_48;
  reg [31:0] GEN_49;
  wire [63:0] T_1198_T_1203_data;
  wire [8:0] T_1198_T_1203_addr;
  wire  T_1198_T_1203_mask;
  wire  T_1198_T_1203_en;
  wire  T_1201;
  wire [8:0] T_1202;
  wire [63:0] GEN_42;
  wire [8:0] T_1204;
  wire [8:0] T_1209;
  reg [63:0] T_1213 [0:511];
  reg [63:0] GEN_50;
  wire [63:0] T_1213_T_1225_data;
  wire [8:0] T_1213_T_1225_addr;
  wire  T_1213_T_1225_en;
  reg [8:0] GEN_51;
  reg [31:0] GEN_52;
  reg  GEN_53;
  reg [31:0] GEN_54;
  wire [63:0] T_1213_T_1218_data;
  wire [8:0] T_1213_T_1218_addr;
  wire  T_1213_T_1218_mask;
  wire  T_1213_T_1218_en;
  wire  T_1216;
  wire [8:0] T_1224;
  reg [63:0] T_1228 [0:511];
  reg [63:0] GEN_55;
  wire [63:0] T_1228_T_1240_data;
  wire [8:0] T_1228_T_1240_addr;
  wire  T_1228_T_1240_en;
  reg [8:0] GEN_56;
  reg [31:0] GEN_57;
  reg  GEN_58;
  reg [31:0] GEN_59;
  wire [63:0] T_1228_T_1233_data;
  wire [8:0] T_1228_T_1233_addr;
  wire  T_1228_T_1233_mask;
  wire  T_1228_T_1233_en;
  wire  T_1231;
  wire [8:0] T_1239;
  reg [63:0] T_1243 [0:511];
  reg [63:0] GEN_60;
  wire [63:0] T_1243_T_1255_data;
  wire [8:0] T_1243_T_1255_addr;
  wire  T_1243_T_1255_en;
  reg [8:0] GEN_61;
  reg [31:0] GEN_62;
  reg  GEN_78;
  reg [31:0] GEN_79;
  wire [63:0] T_1243_T_1248_data;
  wire [8:0] T_1243_T_1248_addr;
  wire  T_1243_T_1248_mask;
  wire  T_1243_T_1248_en;
  wire  T_1246;
  wire [8:0] T_1254;
  wire [63:0] T_1257;
  wire [63:0] T_1259;
  wire [63:0] T_1261;
  wire [63:0] T_1263;
  wire [63:0] T_1265;
  wire [63:0] T_1266;
  wire [63:0] T_1267;
  wire [63:0] T_1268;
  wire  T_1269;
  wire [25:0] T_1270;
  wire [25:0] T_1379_addr_block;
  wire [1:0] T_1379_client_xact_id;
  wire [2:0] T_1379_addr_beat;
  wire  T_1379_is_builtin_type;
  wire [2:0] T_1379_a_type;
  wire [11:0] T_1379_union;
  wire [63:0] T_1379_data;
  wire  T_1410;
  wire [1:0] GEN_63;
  wire [1:0] GEN_64;
  wire  GEN_65;
  wire  T_1412;
  wire [1:0] GEN_66;
  wire [1:0] GEN_67;
  wire  T_1413;
  wire [1:0] GEN_68;
  wire [1:0] GEN_69;
  wire  T_1414;
  wire [1:0] GEN_70;
  wire [1:0] GEN_71;
  reg [31:0] GEN_4;
  reg [31:0] GEN_81;
  FlowThroughSerializer FlowThroughSerializer_1 (
    .clk(FlowThroughSerializer_1_clk),
    .reset(FlowThroughSerializer_1_reset),
    .io_in_ready(FlowThroughSerializer_1_io_in_ready),
    .io_in_valid(FlowThroughSerializer_1_io_in_valid),
    .io_in_bits_addr_beat(FlowThroughSerializer_1_io_in_bits_addr_beat),
    .io_in_bits_client_xact_id(FlowThroughSerializer_1_io_in_bits_client_xact_id),
    .io_in_bits_manager_xact_id(FlowThroughSerializer_1_io_in_bits_manager_xact_id),
    .io_in_bits_is_builtin_type(FlowThroughSerializer_1_io_in_bits_is_builtin_type),
    .io_in_bits_g_type(FlowThroughSerializer_1_io_in_bits_g_type),
    .io_in_bits_data(FlowThroughSerializer_1_io_in_bits_data),
    .io_out_ready(FlowThroughSerializer_1_io_out_ready),
    .io_out_valid(FlowThroughSerializer_1_io_out_valid),
    .io_out_bits_addr_beat(FlowThroughSerializer_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(FlowThroughSerializer_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(FlowThroughSerializer_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(FlowThroughSerializer_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(FlowThroughSerializer_1_io_out_bits_g_type),
    .io_out_bits_data(FlowThroughSerializer_1_io_out_bits_data),
    .io_cnt(FlowThroughSerializer_1_io_cnt),
    .io_done(FlowThroughSerializer_1_io_done)
  );
  assign io_resp_valid = s1_hit;
  assign io_resp_bits_data = GEN_4;
  assign io_resp_bits_datablock = T_1268;
  assign io_mem_acquire_valid = T_1269;
  assign io_mem_acquire_bits_addr_block = T_1379_addr_block;
  assign io_mem_acquire_bits_client_xact_id = T_1379_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = T_1379_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = T_1379_is_builtin_type;
  assign io_mem_acquire_bits_a_type = T_1379_a_type;
  assign io_mem_acquire_bits_union = T_1379_union;
  assign io_mem_acquire_bits_data = T_1379_data;
  assign io_mem_grant_ready = FlowThroughSerializer_1_io_in_ready;
  assign stall = io_resp_ready == 1'h0;
  assign rdy = T_953;
  assign s1_any_tag_hit = T_1195;
  assign T_934 = s1_vaddr[11:0];
  assign s1_paddr = {io_s1_ppn,T_934};
  assign s1_tag = s1_paddr[31:12];
  assign T_935 = s1_valid & stall;
  assign s0_vaddr = T_935 ? s1_vaddr : io_req_bits_addr;
  assign T_937 = io_req_valid & rdy;
  assign T_940 = io_s1_kill == 1'h0;
  assign T_941 = T_935 & T_940;
  assign T_942 = T_937 | T_941;
  assign GEN_0 = T_937 ? io_req_bits_addr : s1_vaddr;
  assign T_946 = s1_valid & T_940;
  assign T_947 = state == 2'h0;
  assign out_valid = T_946 & T_947;
  assign s1_idx = s1_vaddr[11:6];
  assign s1_hit = out_valid & s1_any_tag_hit;
  assign T_949 = s1_any_tag_hit == 1'h0;
  assign s1_miss = out_valid & T_949;
  assign T_952 = s1_miss == 1'h0;
  assign T_953 = T_947 & T_952;
  assign T_955 = s1_valid & T_947;
  assign T_956 = T_955 & s1_miss;
  assign GEN_1 = T_956 ? s1_paddr : refill_addr;
  assign refill_tag = refill_addr[31:12];
  assign FlowThroughSerializer_1_clk = clk;
  assign FlowThroughSerializer_1_reset = reset;
  assign FlowThroughSerializer_1_io_in_valid = io_mem_grant_valid;
  assign FlowThroughSerializer_1_io_in_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign FlowThroughSerializer_1_io_in_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign FlowThroughSerializer_1_io_in_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign FlowThroughSerializer_1_io_in_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign FlowThroughSerializer_1_io_in_bits_g_type = io_mem_grant_bits_g_type;
  assign FlowThroughSerializer_1_io_in_bits_data = io_mem_grant_bits_data;
  assign FlowThroughSerializer_1_io_out_ready = 1'h1;
  assign T_957 = FlowThroughSerializer_1_io_out_ready & FlowThroughSerializer_1_io_out_valid;
  assign T_960 = refill_cnt == 3'h7;
  assign GEN_72 = {{2'd0}, 1'h1};
  assign T_962 = refill_cnt + GEN_72;
  assign T_963 = T_962[2:0];
  assign GEN_2 = T_957 ? T_963 : refill_cnt;
  assign refill_wrap = T_957 & T_960;
  assign T_964 = state == 2'h3;
  assign refill_done = T_964 & refill_wrap;
  assign T_968 = T_967[0];
  assign T_969 = T_967[2];
  assign T_970 = T_968 ^ T_969;
  assign T_971 = T_967[3];
  assign T_972 = T_970 ^ T_971;
  assign T_973 = T_967[5];
  assign T_974 = T_972 ^ T_973;
  assign T_975 = T_967[15:1];
  assign T_976 = {T_974,T_975};
  assign GEN_3 = s1_miss ? T_976 : T_967;
  assign repl_way = T_967[1:0];
  assign tag_array_0_tag_rdata_addr = T_990;
  assign tag_array_0_tag_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_array_0_tag_rdata_data = tag_array_0[GEN_13];
  `else
  assign tag_array_0_tag_rdata_data = GEN_13 >= 7'h40 ? $random : tag_array_0[GEN_13];
  `endif
  assign tag_array_0_T_1018_data = T_999_0;
  assign tag_array_0_T_1018_addr = s1_idx;
  assign tag_array_0_T_1018_mask = GEN_25;
  assign tag_array_0_T_1018_en = refill_done;
  assign tag_array_1_tag_rdata_addr = T_990;
  assign tag_array_1_tag_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_array_1_tag_rdata_data = tag_array_1[GEN_18];
  `else
  assign tag_array_1_tag_rdata_data = GEN_18 >= 7'h40 ? $random : tag_array_1[GEN_18];
  `endif
  assign tag_array_1_T_1018_data = T_999_1;
  assign tag_array_1_T_1018_addr = s1_idx;
  assign tag_array_1_T_1018_mask = GEN_27;
  assign tag_array_1_T_1018_en = refill_done;
  assign tag_array_2_tag_rdata_addr = T_990;
  assign tag_array_2_tag_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_array_2_tag_rdata_data = tag_array_2[GEN_23];
  `else
  assign tag_array_2_tag_rdata_data = GEN_23 >= 7'h40 ? $random : tag_array_2[GEN_23];
  `endif
  assign tag_array_2_T_1018_data = T_999_2;
  assign tag_array_2_T_1018_addr = s1_idx;
  assign tag_array_2_T_1018_mask = GEN_29;
  assign tag_array_2_T_1018_en = refill_done;
  assign tag_array_3_tag_rdata_addr = T_990;
  assign tag_array_3_tag_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_array_3_tag_rdata_data = tag_array_3[GEN_39];
  `else
  assign tag_array_3_tag_rdata_data = GEN_39 >= 7'h40 ? $random : tag_array_3[GEN_39];
  `endif
  assign tag_array_3_T_1018_data = T_999_3;
  assign tag_array_3_T_1018_addr = s1_idx;
  assign tag_array_3_T_1018_mask = GEN_31;
  assign tag_array_3_T_1018_en = refill_done;
  assign T_985 = s0_vaddr[11:6];
  assign T_990 = T_985;
  assign T_999_0 = refill_tag;
  assign T_999_1 = refill_tag;
  assign T_999_2 = refill_tag;
  assign T_999_3 = refill_tag;
  assign GEN_73 = {{1'd0}, 1'h0};
  assign T_1002 = repl_way == GEN_73;
  assign GEN_74 = {{1'd0}, 1'h1};
  assign T_1004 = repl_way == GEN_74;
  assign T_1006 = repl_way == 2'h2;
  assign T_1008 = repl_way == 2'h3;
  assign T_1014_0 = T_1002;
  assign T_1014_1 = T_1004;
  assign T_1014_2 = T_1006;
  assign T_1014_3 = T_1008;
  assign GEN_25 = refill_done ? T_1014_0 : 1'h0;
  assign GEN_27 = refill_done ? T_1014_1 : 1'h0;
  assign GEN_29 = refill_done ? T_1014_2 : 1'h0;
  assign GEN_31 = refill_done ? T_1014_3 : 1'h0;
  assign T_1022 = invalidated == 1'h0;
  assign T_1023 = refill_done & T_1022;
  assign T_1024 = {repl_way,s1_idx};
  assign GEN_75 = {{255'd0}, 1'h1};
  assign T_1027 = GEN_75 << T_1024;
  assign T_1028 = vb_array | T_1027;
  assign T_1029 = ~ vb_array;
  assign GEN_32 = T_1023 ? T_1028 : vb_array;
  assign GEN_33 = io_invalidate ? {{255'd0}, 1'h0} : GEN_32;
  assign GEN_34 = io_invalidate ? 1'h1 : invalidated;
  assign s1_disparity_0 = 1'h0;
  assign s1_disparity_1 = 1'h0;
  assign s1_disparity_2 = 1'h0;
  assign s1_disparity_3 = 1'h0;
  assign T_1042 = s1_valid & s1_disparity_0;
  assign T_1044 = {1'h0,s1_idx};
  assign GEN_76 = {{127'd0}, 1'h1};
  assign T_1047 = GEN_76 << T_1044;
  assign GEN_77 = {{128'd0}, T_1047};
  assign T_1050 = T_1029 | GEN_77;
  assign T_1051 = ~ T_1050;
  assign GEN_35 = T_1042 ? T_1051 : GEN_33;
  assign T_1053 = s1_valid & s1_disparity_1;
  assign T_1055 = {1'h1,s1_idx};
  assign T_1058 = GEN_76 << T_1055;
  assign GEN_80 = {{128'd0}, T_1058};
  assign T_1061 = T_1029 | GEN_80;
  assign T_1062 = ~ T_1061;
  assign GEN_36 = T_1053 ? T_1062 : GEN_35;
  assign T_1064 = s1_valid & s1_disparity_2;
  assign T_1066 = {2'h2,s1_idx};
  assign T_1069 = GEN_75 << T_1066;
  assign T_1072 = T_1029 | T_1069;
  assign T_1073 = ~ T_1072;
  assign GEN_37 = T_1064 ? T_1073 : GEN_36;
  assign T_1075 = s1_valid & s1_disparity_3;
  assign T_1077 = {2'h3,s1_idx};
  assign T_1080 = GEN_75 << T_1077;
  assign T_1083 = T_1029 | T_1080;
  assign T_1084 = ~ T_1083;
  assign GEN_38 = T_1075 ? T_1084 : GEN_37;
  assign s1_tag_match_0 = T_1120;
  assign s1_tag_match_1 = T_1140;
  assign s1_tag_match_2 = T_1160;
  assign s1_tag_match_3 = T_1180;
  assign s1_tag_hit_0 = T_1121;
  assign s1_tag_hit_1 = T_1141;
  assign s1_tag_hit_2 = T_1161;
  assign s1_tag_hit_3 = T_1181;
  assign s1_dout_0 = T_1198_T_1210_data;
  assign s1_dout_1 = T_1213_T_1225_data;
  assign s1_dout_2 = T_1228_T_1240_data;
  assign s1_dout_3 = T_1243_T_1255_data;
  assign T_1108 = io_invalidate == 1'h0;
  assign T_1112 = vb_array >> T_1044;
  assign T_1113 = T_1112[0];
  assign T_1115 = T_1108 & T_1113;
  assign T_1119 = tag_array_0_tag_rdata_data;
  assign T_1120 = T_1119 == s1_tag;
  assign T_1121 = T_1115 & s1_tag_match_0;
  assign T_1132 = vb_array >> T_1055;
  assign T_1133 = T_1132[0];
  assign T_1135 = T_1108 & T_1133;
  assign T_1139 = tag_array_1_tag_rdata_data;
  assign T_1140 = T_1139 == s1_tag;
  assign T_1141 = T_1135 & s1_tag_match_1;
  assign T_1152 = vb_array >> T_1066;
  assign T_1153 = T_1152[0];
  assign T_1155 = T_1108 & T_1153;
  assign T_1159 = tag_array_2_tag_rdata_data;
  assign T_1160 = T_1159 == s1_tag;
  assign T_1161 = T_1155 & s1_tag_match_2;
  assign T_1172 = vb_array >> T_1077;
  assign T_1173 = T_1172[0];
  assign T_1175 = T_1108 & T_1173;
  assign T_1179 = tag_array_3_tag_rdata_data;
  assign T_1180 = T_1179 == s1_tag;
  assign T_1181 = T_1175 & s1_tag_match_3;
  assign T_1187 = s1_tag_hit_0 | s1_tag_hit_1;
  assign T_1188 = T_1187 | s1_tag_hit_2;
  assign T_1189 = T_1188 | s1_tag_hit_3;
  assign T_1190 = s1_disparity_0 | s1_disparity_1;
  assign T_1191 = T_1190 | s1_disparity_2;
  assign T_1192 = T_1191 | s1_disparity_3;
  assign T_1194 = T_1192 == 1'h0;
  assign T_1195 = T_1189 & T_1194;
  assign T_1198_T_1210_addr = T_1209;
  assign T_1198_T_1210_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1198_T_1210_data = T_1198[GEN_46];
  `else
  assign T_1198_T_1210_data = GEN_46 >= 10'h200 ? $random : T_1198[GEN_46];
  `endif
  assign T_1198_T_1203_data = GEN_42;
  assign T_1198_T_1203_addr = T_1202;
  assign T_1198_T_1203_mask = T_1201;
  assign T_1198_T_1203_en = T_1201;
  assign T_1201 = FlowThroughSerializer_1_io_out_valid & T_1002;
  assign T_1202 = {s1_idx,refill_cnt};
  assign GEN_42 = FlowThroughSerializer_1_io_out_bits_data;
  assign T_1204 = s0_vaddr[11:3];
  assign T_1209 = T_1204;
  assign T_1213_T_1225_addr = T_1224;
  assign T_1213_T_1225_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1213_T_1225_data = T_1213[GEN_51];
  `else
  assign T_1213_T_1225_data = GEN_51 >= 10'h200 ? $random : T_1213[GEN_51];
  `endif
  assign T_1213_T_1218_data = GEN_42;
  assign T_1213_T_1218_addr = T_1202;
  assign T_1213_T_1218_mask = T_1216;
  assign T_1213_T_1218_en = T_1216;
  assign T_1216 = FlowThroughSerializer_1_io_out_valid & T_1004;
  assign T_1224 = T_1204;
  assign T_1228_T_1240_addr = T_1239;
  assign T_1228_T_1240_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1228_T_1240_data = T_1228[GEN_56];
  `else
  assign T_1228_T_1240_data = GEN_56 >= 10'h200 ? $random : T_1228[GEN_56];
  `endif
  assign T_1228_T_1233_data = GEN_42;
  assign T_1228_T_1233_addr = T_1202;
  assign T_1228_T_1233_mask = T_1231;
  assign T_1228_T_1233_en = T_1231;
  assign T_1231 = FlowThroughSerializer_1_io_out_valid & T_1006;
  assign T_1239 = T_1204;
  assign T_1243_T_1255_addr = T_1254;
  assign T_1243_T_1255_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1243_T_1255_data = T_1243[GEN_61];
  `else
  assign T_1243_T_1255_data = GEN_61 >= 10'h200 ? $random : T_1243[GEN_61];
  `endif
  assign T_1243_T_1248_data = GEN_42;
  assign T_1243_T_1248_addr = T_1202;
  assign T_1243_T_1248_mask = T_1246;
  assign T_1243_T_1248_en = T_1246;
  assign T_1246 = FlowThroughSerializer_1_io_out_valid & T_1008;
  assign T_1254 = T_1204;
  assign T_1257 = s1_tag_hit_0 ? s1_dout_0 : {{63'd0}, 1'h0};
  assign T_1259 = s1_tag_hit_1 ? s1_dout_1 : {{63'd0}, 1'h0};
  assign T_1261 = s1_tag_hit_2 ? s1_dout_2 : {{63'd0}, 1'h0};
  assign T_1263 = s1_tag_hit_3 ? s1_dout_3 : {{63'd0}, 1'h0};
  assign T_1265 = T_1257 | T_1259;
  assign T_1266 = T_1265 | T_1261;
  assign T_1267 = T_1266 | T_1263;
  assign T_1268 = T_1267;
  assign T_1269 = state == 2'h1;
  assign T_1270 = refill_addr[31:6];
  assign T_1379_addr_block = T_1270;
  assign T_1379_client_xact_id = {{1'd0}, 1'h0};
  assign T_1379_addr_beat = {{2'd0}, 1'h0};
  assign T_1379_is_builtin_type = 1'h1;
  assign T_1379_a_type = 3'h1;
  assign T_1379_union = 12'h1c1;
  assign T_1379_data = {{63'd0}, 1'h0};
  assign T_1410 = 2'h0 == state;
  assign GEN_63 = s1_miss ? 2'h1 : state;
  assign GEN_64 = T_1410 ? GEN_63 : state;
  assign GEN_65 = T_1410 ? 1'h0 : GEN_34;
  assign T_1412 = 2'h1 == state;
  assign GEN_66 = io_mem_acquire_ready ? 2'h2 : GEN_64;
  assign GEN_67 = T_1412 ? GEN_66 : GEN_64;
  assign T_1413 = 2'h2 == state;
  assign GEN_68 = io_mem_grant_valid ? 2'h3 : GEN_67;
  assign GEN_69 = T_1413 ? GEN_68 : GEN_67;
  assign T_1414 = 2'h3 == state;
  assign GEN_70 = refill_done ? 2'h0 : GEN_69;
  assign GEN_71 = T_1414 ? GEN_70 : GEN_69;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_5 = {1{$random}};
  state = GEN_5[1:0];
  GEN_6 = {1{$random}};
  invalidated = GEN_6[0:0];
  GEN_7 = {1{$random}};
  refill_addr = GEN_7[31:0];
  GEN_8 = {1{$random}};
  s1_valid = GEN_8[0:0];
  GEN_9 = {2{$random}};
  s1_vaddr = GEN_9[38:0];
  GEN_10 = {1{$random}};
  refill_cnt = GEN_10[2:0];
  GEN_11 = {1{$random}};
  T_967 = GEN_11[15:0];
  GEN_12 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = GEN_12[19:0];
  GEN_14 = {1{$random}};
  GEN_13 = GEN_14[5:0];
  GEN_16 = {1{$random}};
  GEN_15 = GEN_16[0:0];
  GEN_17 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = GEN_17[19:0];
  GEN_19 = {1{$random}};
  GEN_18 = GEN_19[5:0];
  GEN_21 = {1{$random}};
  GEN_20 = GEN_21[0:0];
  GEN_22 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = GEN_22[19:0];
  GEN_24 = {1{$random}};
  GEN_23 = GEN_24[5:0];
  GEN_28 = {1{$random}};
  GEN_26 = GEN_28[0:0];
  GEN_30 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = GEN_30[19:0];
  GEN_40 = {1{$random}};
  GEN_39 = GEN_40[5:0];
  GEN_43 = {1{$random}};
  GEN_41 = GEN_43[0:0];
  GEN_44 = {8{$random}};
  vb_array = GEN_44[255:0];
  GEN_45 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1198[initvar] = GEN_45[63:0];
  GEN_47 = {1{$random}};
  GEN_46 = GEN_47[8:0];
  GEN_49 = {1{$random}};
  GEN_48 = GEN_49[0:0];
  GEN_50 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1213[initvar] = GEN_50[63:0];
  GEN_52 = {1{$random}};
  GEN_51 = GEN_52[8:0];
  GEN_54 = {1{$random}};
  GEN_53 = GEN_54[0:0];
  GEN_55 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1228[initvar] = GEN_55[63:0];
  GEN_57 = {1{$random}};
  GEN_56 = GEN_57[8:0];
  GEN_59 = {1{$random}};
  GEN_58 = GEN_59[0:0];
  GEN_60 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1243[initvar] = GEN_60[63:0];
  GEN_62 = {1{$random}};
  GEN_61 = GEN_62[8:0];
  GEN_79 = {1{$random}};
  GEN_78 = GEN_79[0:0];
  GEN_81 = {1{$random}};
  GEN_4 = GEN_81[31:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else begin
      if(T_1414) begin
        if(refill_done) begin
          state <= 2'h0;
        end else begin
          if(T_1413) begin
            if(io_mem_grant_valid) begin
              state <= 2'h3;
            end else begin
              if(T_1412) begin
                if(io_mem_acquire_ready) begin
                  state <= 2'h2;
                end else begin
                  if(T_1410) begin
                    if(s1_miss) begin
                      state <= 2'h1;
                    end
                  end
                end
              end else begin
                if(T_1410) begin
                  if(s1_miss) begin
                    state <= 2'h1;
                  end
                end
              end
            end
          end else begin
            if(T_1412) begin
              if(io_mem_acquire_ready) begin
                state <= 2'h2;
              end else begin
                if(T_1410) begin
                  if(s1_miss) begin
                    state <= 2'h1;
                  end
                end
              end
            end else begin
              if(T_1410) begin
                if(s1_miss) begin
                  state <= 2'h1;
                end
              end
            end
          end
        end
      end else begin
        if(T_1413) begin
          if(io_mem_grant_valid) begin
            state <= 2'h3;
          end else begin
            if(T_1412) begin
              if(io_mem_acquire_ready) begin
                state <= 2'h2;
              end else begin
                state <= GEN_64;
              end
            end else begin
              state <= GEN_64;
            end
          end
        end else begin
          if(T_1412) begin
            if(io_mem_acquire_ready) begin
              state <= 2'h2;
            end else begin
              state <= GEN_64;
            end
          end else begin
            state <= GEN_64;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1410) begin
        invalidated <= 1'h0;
      end else begin
        if(io_invalidate) begin
          invalidated <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_956) begin
        refill_addr <= s1_paddr;
      end
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_942;
    end
    if(1'h0) begin
    end else begin
      if(T_937) begin
        s1_vaddr <= io_req_bits_addr;
      end
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      if(T_957) begin
        refill_cnt <= T_963;
      end
    end
    if(reset) begin
      T_967 <= 16'h1;
    end else begin
      if(s1_miss) begin
        T_967 <= T_976;
      end
    end
    GEN_13 <= tag_array_0_tag_rdata_addr;
    GEN_15 <= tag_array_0_tag_rdata_en;
    if(tag_array_0_T_1018_en & tag_array_0_T_1018_mask) begin
      tag_array_0[tag_array_0_T_1018_addr] <= tag_array_0_T_1018_data;
    end
    GEN_18 <= tag_array_1_tag_rdata_addr;
    GEN_20 <= tag_array_1_tag_rdata_en;
    if(tag_array_1_T_1018_en & tag_array_1_T_1018_mask) begin
      tag_array_1[tag_array_1_T_1018_addr] <= tag_array_1_T_1018_data;
    end
    GEN_23 <= tag_array_2_tag_rdata_addr;
    GEN_26 <= tag_array_2_tag_rdata_en;
    if(tag_array_2_T_1018_en & tag_array_2_T_1018_mask) begin
      tag_array_2[tag_array_2_T_1018_addr] <= tag_array_2_T_1018_data;
    end
    GEN_39 <= tag_array_3_tag_rdata_addr;
    GEN_41 <= tag_array_3_tag_rdata_en;
    if(tag_array_3_T_1018_en & tag_array_3_T_1018_mask) begin
      tag_array_3[tag_array_3_T_1018_addr] <= tag_array_3_T_1018_data;
    end
    if(reset) begin
      vb_array <= 256'h0;
    end else begin
      if(T_1075) begin
        vb_array <= T_1084;
      end else begin
        if(T_1064) begin
          vb_array <= T_1073;
        end else begin
          if(T_1053) begin
            vb_array <= T_1062;
          end else begin
            if(T_1042) begin
              vb_array <= T_1051;
            end else begin
              if(io_invalidate) begin
                vb_array <= {{255'd0}, 1'h0};
              end else begin
                if(T_1023) begin
                  vb_array <= T_1028;
                end
              end
            end
          end
        end
      end
    end
    GEN_46 <= T_1198_T_1210_addr;
    GEN_48 <= T_1198_T_1210_en;
    if(T_1198_T_1203_en & T_1198_T_1203_mask) begin
      T_1198[T_1198_T_1203_addr] <= T_1198_T_1203_data;
    end
    GEN_51 <= T_1213_T_1225_addr;
    GEN_53 <= T_1213_T_1225_en;
    if(T_1213_T_1218_en & T_1213_T_1218_mask) begin
      T_1213[T_1213_T_1218_addr] <= T_1213_T_1218_data;
    end
    GEN_56 <= T_1228_T_1240_addr;
    GEN_58 <= T_1228_T_1240_en;
    if(T_1228_T_1233_en & T_1228_T_1233_mask) begin
      T_1228[T_1228_T_1233_addr] <= T_1228_T_1233_data;
    end
    GEN_61 <= T_1243_T_1255_addr;
    GEN_78 <= T_1243_T_1255_en;
    if(T_1243_T_1248_en & T_1243_T_1248_mask) begin
      T_1243[T_1243_T_1248_addr] <= T_1243_T_1248_data;
    end
  end
endmodule
module RocketCAM(
  input   clk,
  input   reset,
  input   io_clear,
  input  [7:0] io_clear_mask,
  input  [33:0] io_tag,
  output  io_hit,
  output [7:0] io_hits,
  output [7:0] io_valid_bits,
  input   io_write,
  input  [33:0] io_write_tag,
  input  [2:0] io_write_addr
);
  reg [33:0] cam_tags [0:7];
  reg [63:0] GEN_1;
  wire [33:0] cam_tags_T_25_data;
  wire [2:0] cam_tags_T_25_addr;
  wire  cam_tags_T_25_en;
  wire [33:0] cam_tags_T_30_data;
  wire [2:0] cam_tags_T_30_addr;
  wire  cam_tags_T_30_en;
  wire [33:0] cam_tags_T_35_data;
  wire [2:0] cam_tags_T_35_addr;
  wire  cam_tags_T_35_en;
  wire [33:0] cam_tags_T_40_data;
  wire [2:0] cam_tags_T_40_addr;
  wire  cam_tags_T_40_en;
  wire [33:0] cam_tags_T_45_data;
  wire [2:0] cam_tags_T_45_addr;
  wire  cam_tags_T_45_en;
  wire [33:0] cam_tags_T_50_data;
  wire [2:0] cam_tags_T_50_addr;
  wire  cam_tags_T_50_en;
  wire [33:0] cam_tags_T_55_data;
  wire [2:0] cam_tags_T_55_addr;
  wire  cam_tags_T_55_en;
  wire [33:0] cam_tags_T_60_data;
  wire [2:0] cam_tags_T_60_addr;
  wire  cam_tags_T_60_en;
  wire [33:0] cam_tags_T_20_data;
  wire [2:0] cam_tags_T_20_addr;
  wire  cam_tags_T_20_mask;
  wire  cam_tags_T_20_en;
  reg [7:0] vb_array;
  reg [31:0] GEN_2;
  wire [7:0] GEN_7;
  wire [7:0] T_14;
  wire [7:0] T_15;
  wire [7:0] GEN_0;
  wire [7:0] T_21;
  wire [7:0] T_22;
  wire [7:0] GEN_6;
  wire  T_23;
  wire  T_26;
  wire  T_27;
  wire  T_28;
  wire  T_31;
  wire  T_32;
  wire  T_33;
  wire  T_36;
  wire  T_37;
  wire  T_38;
  wire  T_41;
  wire  T_42;
  wire  T_43;
  wire  T_46;
  wire  T_47;
  wire  T_48;
  wire  T_51;
  wire  T_52;
  wire  T_53;
  wire  T_56;
  wire  T_57;
  wire  T_58;
  wire  T_61;
  wire  T_62;
  wire  T_68_0;
  wire  T_68_1;
  wire  T_68_2;
  wire  T_68_3;
  wire  T_68_4;
  wire  T_68_5;
  wire  T_68_6;
  wire  T_68_7;
  wire [1:0] T_70;
  wire [1:0] T_71;
  wire [3:0] T_72;
  wire [1:0] T_73;
  wire [1:0] T_74;
  wire [3:0] T_75;
  wire [7:0] T_76;
  wire [7:0] GEN_8;
  wire  T_78;
  assign io_hit = T_78;
  assign io_hits = T_76;
  assign io_valid_bits = vb_array;
  assign cam_tags_T_25_addr = {{2'd0}, 1'h0};
  assign cam_tags_T_25_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_25_data = cam_tags[cam_tags_T_25_addr];
  `else
  assign cam_tags_T_25_data = cam_tags_T_25_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_25_addr];
  `endif
  assign cam_tags_T_30_addr = {{2'd0}, 1'h1};
  assign cam_tags_T_30_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_30_data = cam_tags[cam_tags_T_30_addr];
  `else
  assign cam_tags_T_30_data = cam_tags_T_30_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_30_addr];
  `endif
  assign cam_tags_T_35_addr = {{1'd0}, 2'h2};
  assign cam_tags_T_35_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_35_data = cam_tags[cam_tags_T_35_addr];
  `else
  assign cam_tags_T_35_data = cam_tags_T_35_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_35_addr];
  `endif
  assign cam_tags_T_40_addr = {{1'd0}, 2'h3};
  assign cam_tags_T_40_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_40_data = cam_tags[cam_tags_T_40_addr];
  `else
  assign cam_tags_T_40_data = cam_tags_T_40_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_40_addr];
  `endif
  assign cam_tags_T_45_addr = 3'h4;
  assign cam_tags_T_45_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_45_data = cam_tags[cam_tags_T_45_addr];
  `else
  assign cam_tags_T_45_data = cam_tags_T_45_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_45_addr];
  `endif
  assign cam_tags_T_50_addr = 3'h5;
  assign cam_tags_T_50_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_50_data = cam_tags[cam_tags_T_50_addr];
  `else
  assign cam_tags_T_50_data = cam_tags_T_50_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_50_addr];
  `endif
  assign cam_tags_T_55_addr = 3'h6;
  assign cam_tags_T_55_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_55_data = cam_tags[cam_tags_T_55_addr];
  `else
  assign cam_tags_T_55_data = cam_tags_T_55_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_55_addr];
  `endif
  assign cam_tags_T_60_addr = 3'h7;
  assign cam_tags_T_60_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_60_data = cam_tags[cam_tags_T_60_addr];
  `else
  assign cam_tags_T_60_data = cam_tags_T_60_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_60_addr];
  `endif
  assign cam_tags_T_20_data = io_write_tag;
  assign cam_tags_T_20_addr = io_write_addr;
  assign cam_tags_T_20_mask = io_write;
  assign cam_tags_T_20_en = io_write;
  assign GEN_7 = {{7'd0}, 1'h1};
  assign T_14 = GEN_7 << io_write_addr;
  assign T_15 = vb_array | T_14;
  assign GEN_0 = io_write ? T_15 : vb_array;
  assign T_21 = ~ io_clear_mask;
  assign T_22 = vb_array & T_21;
  assign GEN_6 = io_clear ? T_22 : GEN_0;
  assign T_23 = vb_array[0];
  assign T_26 = cam_tags_T_25_data == io_tag;
  assign T_27 = T_23 & T_26;
  assign T_28 = vb_array[1];
  assign T_31 = cam_tags_T_30_data == io_tag;
  assign T_32 = T_28 & T_31;
  assign T_33 = vb_array[2];
  assign T_36 = cam_tags_T_35_data == io_tag;
  assign T_37 = T_33 & T_36;
  assign T_38 = vb_array[3];
  assign T_41 = cam_tags_T_40_data == io_tag;
  assign T_42 = T_38 & T_41;
  assign T_43 = vb_array[4];
  assign T_46 = cam_tags_T_45_data == io_tag;
  assign T_47 = T_43 & T_46;
  assign T_48 = vb_array[5];
  assign T_51 = cam_tags_T_50_data == io_tag;
  assign T_52 = T_48 & T_51;
  assign T_53 = vb_array[6];
  assign T_56 = cam_tags_T_55_data == io_tag;
  assign T_57 = T_53 & T_56;
  assign T_58 = vb_array[7];
  assign T_61 = cam_tags_T_60_data == io_tag;
  assign T_62 = T_58 & T_61;
  assign T_68_0 = T_27;
  assign T_68_1 = T_32;
  assign T_68_2 = T_37;
  assign T_68_3 = T_42;
  assign T_68_4 = T_47;
  assign T_68_5 = T_52;
  assign T_68_6 = T_57;
  assign T_68_7 = T_62;
  assign T_70 = {T_68_1,T_68_0};
  assign T_71 = {T_68_3,T_68_2};
  assign T_72 = {T_71,T_70};
  assign T_73 = {T_68_5,T_68_4};
  assign T_74 = {T_68_7,T_68_6};
  assign T_75 = {T_74,T_73};
  assign T_76 = {T_75,T_72};
  assign GEN_8 = {{7'd0}, 1'h0};
  assign T_78 = io_hits != GEN_8;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_1 = {2{$random}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cam_tags[initvar] = GEN_1[33:0];
  GEN_2 = {1{$random}};
  vb_array = GEN_2[7:0];
  end
`endif
  always @(posedge clk) begin
    if(cam_tags_T_20_en & cam_tags_T_20_mask) begin
      cam_tags[cam_tags_T_20_addr] <= cam_tags_T_20_data;
    end
    if(reset) begin
      vb_array <= 8'h0;
    end else begin
      if(io_clear) begin
        vb_array <= T_22;
      end else begin
        if(io_write) begin
          vb_array <= T_15;
        end
      end
    end
  end
endmodule
module TLB(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [27:0] io_req_bits_vpn,
  input   io_req_bits_passthrough,
  input   io_req_bits_instruction,
  input   io_req_bits_store,
  output  io_resp_miss,
  output [19:0] io_resp_ppn,
  output  io_resp_xcpt_ld,
  output  io_resp_xcpt_st,
  output  io_resp_xcpt_if,
  output [7:0] io_resp_hit_idx,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_addr,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [19:0] io_ptw_resp_bits_pte_ppn,
  input  [2:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_r,
  input  [3:0] io_ptw_resp_bits_pte_typ,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [4:0] io_ptw_status_zero1,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie
);
  wire  tag_cam_clk;
  wire  tag_cam_reset;
  wire  tag_cam_io_clear;
  wire [7:0] tag_cam_io_clear_mask;
  wire [33:0] tag_cam_io_tag;
  wire  tag_cam_io_hit;
  wire [7:0] tag_cam_io_hits;
  wire [7:0] tag_cam_io_valid_bits;
  wire  tag_cam_io_write;
  wire [33:0] tag_cam_io_write_tag;
  wire [2:0] tag_cam_io_write_addr;
  reg [19:0] tag_ram [0:7];
  reg [31:0] GEN_63;
  wire [19:0] tag_ram_T_561_data;
  wire [2:0] tag_ram_T_561_addr;
  wire  tag_ram_T_561_en;
  wire [19:0] tag_ram_T_563_data;
  wire [2:0] tag_ram_T_563_addr;
  wire  tag_ram_T_563_en;
  wire [19:0] tag_ram_T_565_data;
  wire [2:0] tag_ram_T_565_addr;
  wire  tag_ram_T_565_en;
  wire [19:0] tag_ram_T_567_data;
  wire [2:0] tag_ram_T_567_addr;
  wire  tag_ram_T_567_en;
  wire [19:0] tag_ram_T_569_data;
  wire [2:0] tag_ram_T_569_addr;
  wire  tag_ram_T_569_en;
  wire [19:0] tag_ram_T_571_data;
  wire [2:0] tag_ram_T_571_addr;
  wire  tag_ram_T_571_en;
  wire [19:0] tag_ram_T_573_data;
  wire [2:0] tag_ram_T_573_addr;
  wire  tag_ram_T_573_en;
  wire [19:0] tag_ram_T_575_data;
  wire [2:0] tag_ram_T_575_addr;
  wire  tag_ram_T_575_en;
  wire [19:0] tag_ram_T_231_data;
  wire [2:0] tag_ram_T_231_addr;
  wire  tag_ram_T_231_mask;
  wire  tag_ram_T_231_en;
  reg [1:0] state;
  reg [31:0] GEN_64;
  reg [33:0] r_refill_tag;
  reg [63:0] GEN_65;
  reg [2:0] r_refill_waddr;
  reg [31:0] GEN_66;
  reg [27:0] r_req_vpn;
  reg [31:0] GEN_67;
  reg  r_req_passthrough;
  reg [31:0] GEN_68;
  reg  r_req_instruction;
  reg [31:0] GEN_77;
  reg  r_req_store;
  reg [31:0] GEN_86;
  wire [26:0] T_167;
  wire [33:0] lookup_tag;
  wire  T_168;
  wire  T_169;
  wire [3:0] T_170;
  wire [3:0] T_171;
  wire [3:0] GEN_145;
  wire  T_173;
  wire [3:0] T_174;
  wire [1:0] T_175;
  wire [1:0] T_176;
  wire [1:0] GEN_146;
  wire  T_178;
  wire [1:0] T_179;
  wire  T_180;
  wire [1:0] T_181;
  wire [2:0] tag_hit_addr;
  reg  ur_array_0;
  reg [31:0] GEN_95;
  reg  ur_array_1;
  reg [31:0] GEN_104;
  reg  ur_array_2;
  reg [31:0] GEN_113;
  reg  ur_array_3;
  reg [31:0] GEN_122;
  reg  ur_array_4;
  reg [31:0] GEN_152;
  reg  ur_array_5;
  reg [31:0] GEN_153;
  reg  ur_array_6;
  reg [31:0] GEN_154;
  reg  ur_array_7;
  reg [31:0] GEN_155;
  reg  uw_array_0;
  reg [31:0] GEN_156;
  reg  uw_array_1;
  reg [31:0] GEN_157;
  reg  uw_array_2;
  reg [31:0] GEN_158;
  reg  uw_array_3;
  reg [31:0] GEN_159;
  reg  uw_array_4;
  reg [31:0] GEN_160;
  reg  uw_array_5;
  reg [31:0] GEN_161;
  reg  uw_array_6;
  reg [31:0] GEN_162;
  reg  uw_array_7;
  reg [31:0] GEN_163;
  reg  ux_array_0;
  reg [31:0] GEN_164;
  reg  ux_array_1;
  reg [31:0] GEN_165;
  reg  ux_array_2;
  reg [31:0] GEN_166;
  reg  ux_array_3;
  reg [31:0] GEN_167;
  reg  ux_array_4;
  reg [31:0] GEN_168;
  reg  ux_array_5;
  reg [31:0] GEN_169;
  reg  ux_array_6;
  reg [31:0] GEN_170;
  reg  ux_array_7;
  reg [31:0] GEN_171;
  reg  sr_array_0;
  reg [31:0] GEN_173;
  reg  sr_array_1;
  reg [31:0] GEN_174;
  reg  sr_array_2;
  reg [31:0] GEN_175;
  reg  sr_array_3;
  reg [31:0] GEN_176;
  reg  sr_array_4;
  reg [31:0] GEN_177;
  reg  sr_array_5;
  reg [31:0] GEN_178;
  reg  sr_array_6;
  reg [31:0] GEN_179;
  reg  sr_array_7;
  reg [31:0] GEN_180;
  reg  sw_array_0;
  reg [31:0] GEN_183;
  reg  sw_array_1;
  reg [31:0] GEN_184;
  reg  sw_array_2;
  reg [31:0] GEN_185;
  reg  sw_array_3;
  reg [31:0] GEN_186;
  reg  sw_array_4;
  reg [31:0] GEN_191;
  reg  sw_array_5;
  reg [31:0] GEN_193;
  reg  sw_array_6;
  reg [31:0] GEN_197;
  reg  sw_array_7;
  reg [31:0] GEN_200;
  reg  sx_array_0;
  reg [31:0] GEN_201;
  reg  sx_array_1;
  reg [31:0] GEN_202;
  reg  sx_array_2;
  reg [31:0] GEN_203;
  reg  sx_array_3;
  reg [31:0] GEN_204;
  reg  sx_array_4;
  reg [31:0] GEN_205;
  reg  sx_array_5;
  reg [31:0] GEN_206;
  reg  sx_array_6;
  reg [31:0] GEN_207;
  reg  sx_array_7;
  reg [31:0] GEN_208;
  reg  dirty_array_0;
  reg [31:0] GEN_209;
  reg  dirty_array_1;
  reg [31:0] GEN_210;
  reg  dirty_array_2;
  reg [31:0] GEN_211;
  reg  dirty_array_3;
  reg [31:0] GEN_212;
  reg  dirty_array_4;
  reg [31:0] GEN_213;
  reg  dirty_array_5;
  reg [31:0] GEN_214;
  reg  dirty_array_6;
  reg [31:0] GEN_215;
  reg  dirty_array_7;
  reg [31:0] GEN_216;
  wire [3:0] GEN_147;
  wire  T_233;
  wire  T_234;
  wire  T_236;
  wire  T_237;
  wire  GEN_0;
  wire [2:0] GEN_148;
  wire  GEN_7;
  wire [2:0] GEN_149;
  wire  GEN_8;
  wire [2:0] GEN_150;
  wire  GEN_9;
  wire [2:0] GEN_151;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  T_244;
  wire  T_245;
  wire  GEN_1;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  T_252;
  wire  T_253;
  wire  GEN_2;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_3;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  T_261;
  wire  GEN_4;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire [3:0] GEN_172;
  wire  T_263;
  wire  T_264;
  wire  T_266;
  wire  GEN_5;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_6;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire  GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_62;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire [7:0] T_267;
  wire [7:0] GEN_181;
  wire  T_269;
  wire  has_invalid_entry;
  wire  T_272;
  wire  T_273;
  wire  T_274;
  wire  T_275;
  wire  T_276;
  wire  T_277;
  wire  T_278;
  wire [2:0] T_288;
  wire [2:0] T_289;
  wire [2:0] T_290;
  wire [2:0] T_291;
  wire [2:0] T_292;
  wire [2:0] T_293;
  wire [2:0] invalid_entry;
  reg [7:0] T_295;
  reg [31:0] GEN_217;
  wire [7:0] T_297;
  wire  T_298;
  wire [1:0] T_299;
  wire [7:0] T_300;
  wire  T_301;
  wire [2:0] T_302;
  wire [7:0] T_303;
  wire  T_304;
  wire [3:0] T_305;
  wire [2:0] T_306;
  wire [2:0] repl_waddr;
  wire  T_308;
  wire  do_mprv;
  wire [1:0] priv;
  wire [1:0] GEN_182;
  wire  priv_s;
  wire  T_311;
  wire  T_313;
  wire  priv_uses_vm;
  wire [1:0] T_320;
  wire [1:0] T_321;
  wire [3:0] T_322;
  wire [1:0] T_323;
  wire [1:0] T_324;
  wire [3:0] T_325;
  wire [7:0] ur_bits;
  wire [7:0] T_327;
  wire [7:0] pum_ok;
  wire [1:0] T_328;
  wire [1:0] T_329;
  wire [3:0] T_330;
  wire [1:0] T_331;
  wire [1:0] T_332;
  wire [3:0] T_333;
  wire [7:0] T_334;
  wire [7:0] T_335;
  wire [7:0] r_array;
  wire [1:0] T_336;
  wire [1:0] T_337;
  wire [3:0] T_338;
  wire [1:0] T_339;
  wire [1:0] T_340;
  wire [3:0] T_341;
  wire [7:0] T_342;
  wire [7:0] T_343;
  wire [1:0] T_344;
  wire [1:0] T_345;
  wire [3:0] T_346;
  wire [1:0] T_347;
  wire [1:0] T_348;
  wire [3:0] T_349;
  wire [7:0] T_350;
  wire [7:0] w_array;
  wire [1:0] T_351;
  wire [1:0] T_352;
  wire [3:0] T_353;
  wire [1:0] T_354;
  wire [1:0] T_355;
  wire [3:0] T_356;
  wire [7:0] T_357;
  wire [1:0] T_358;
  wire [1:0] T_359;
  wire [3:0] T_360;
  wire [1:0] T_361;
  wire [1:0] T_362;
  wire [3:0] T_363;
  wire [7:0] T_364;
  wire [7:0] x_array;
  wire  T_366;
  wire  T_368;
  wire  T_370;
  wire  vm_enabled;
  wire  T_371;
  wire  T_372;
  wire  bad_va;
  wire [1:0] T_373;
  wire [1:0] T_374;
  wire [3:0] T_375;
  wire [1:0] T_376;
  wire [1:0] T_377;
  wire [3:0] T_378;
  wire [7:0] T_379;
  wire [7:0] T_381;
  wire [7:0] T_382;
  wire [7:0] T_383;
  wire [7:0] tag_hits;
  wire  tag_hit;
  wire  tlb_hit;
  wire  T_386;
  wire  T_387;
  wire  T_389;
  wire  tlb_miss;
  wire  T_390;
  wire  T_405;
  wire [8:0] GEN_187;
  wire [8:0] T_407;
  wire [7:0] T_408;
  wire [7:0] T_409;
  wire [7:0] T_410;
  wire [7:0] T_412;
  wire [7:0] T_413;
  wire [1:0] T_414;
  wire  T_415;
  wire [10:0] GEN_188;
  wire [10:0] T_417;
  wire [7:0] T_418;
  wire [7:0] T_419;
  wire [7:0] T_420;
  wire [7:0] T_422;
  wire [7:0] T_423;
  wire [2:0] T_424;
  wire  T_425;
  wire [14:0] GEN_189;
  wire [14:0] T_427;
  wire [7:0] T_428;
  wire [7:0] T_429;
  wire [7:0] T_430;
  wire [7:0] T_432;
  wire [7:0] T_433;
  wire [7:0] GEN_131;
  wire [31:0] paddr;
  wire [31:0] GEN_190;
  wire  T_439;
  wire [2:0] T_443;
  wire  T_445;
  wire [31:0] GEN_192;
  wire  T_447;
  wire  T_448;
  wire [2:0] T_451;
  wire  T_453;
  wire [31:0] GEN_194;
  wire  T_455;
  wire  T_456;
  wire [2:0] T_459;
  wire [31:0] GEN_195;
  wire  T_461;
  wire [31:0] GEN_196;
  wire  T_463;
  wire  T_464;
  wire [2:0] T_467;
  wire  T_469;
  wire [31:0] GEN_198;
  wire  T_471;
  wire  T_472;
  wire [2:0] T_475;
  wire [31:0] GEN_199;
  wire  T_477;
  wire  T_479;
  wire  T_480;
  wire [2:0] T_483;
  wire  T_485;
  wire [2:0] T_491;
  wire [2:0] T_496;
  wire [2:0] T_497;
  wire [2:0] T_498;
  wire [2:0] T_499;
  wire [2:0] T_500;
  wire [2:0] T_501;
  wire  addr_prot_x;
  wire  addr_prot_w;
  wire  addr_prot_r;
  wire  T_509;
  wire  T_510;
  wire  T_511;
  wire  T_512;
  wire  T_514;
  wire  T_516;
  wire  T_517;
  wire  T_518;
  wire [7:0] T_519;
  wire  T_521;
  wire  T_523;
  wire  T_524;
  wire  T_525;
  wire  T_529;
  wire  T_530;
  wire  T_531;
  wire [7:0] T_532;
  wire  T_534;
  wire  T_536;
  wire  T_537;
  wire  T_538;
  wire  T_542;
  wire  T_543;
  wire  T_544;
  wire [7:0] T_545;
  wire  T_547;
  wire  T_549;
  wire  T_550;
  wire  T_551;
  wire  T_552;
  wire  T_553;
  wire  T_554;
  wire  T_555;
  wire  T_556;
  wire  T_557;
  wire  T_558;
  wire  T_559;
  wire [19:0] T_577;
  wire [19:0] T_579;
  wire [19:0] T_581;
  wire [19:0] T_583;
  wire [19:0] T_585;
  wire [19:0] T_587;
  wire [19:0] T_589;
  wire [19:0] T_591;
  wire [19:0] T_593;
  wire [19:0] T_594;
  wire [19:0] T_595;
  wire [19:0] T_596;
  wire [19:0] T_597;
  wire [19:0] T_598;
  wire [19:0] T_599;
  wire [19:0] T_600;
  wire [19:0] T_601;
  wire [19:0] T_602;
  wire  T_605;
  wire  T_606;
  wire  T_607;
  wire [1:0] GEN_132;
  wire [33:0] GEN_133;
  wire [2:0] GEN_134;
  wire [27:0] GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire [1:0] GEN_139;
  wire [1:0] GEN_140;
  wire [1:0] GEN_141;
  wire [1:0] GEN_142;
  wire  T_610;
  wire [1:0] GEN_143;
  wire [1:0] GEN_144;
  RocketCAM tag_cam (
    .clk(tag_cam_clk),
    .reset(tag_cam_reset),
    .io_clear(tag_cam_io_clear),
    .io_clear_mask(tag_cam_io_clear_mask),
    .io_tag(tag_cam_io_tag),
    .io_hit(tag_cam_io_hit),
    .io_hits(tag_cam_io_hits),
    .io_valid_bits(tag_cam_io_valid_bits),
    .io_write(tag_cam_io_write),
    .io_write_tag(tag_cam_io_write_tag),
    .io_write_addr(tag_cam_io_write_addr)
  );
  assign io_req_ready = T_512;
  assign io_resp_miss = tlb_miss;
  assign io_resp_ppn = T_602;
  assign io_resp_xcpt_ld = T_525;
  assign io_resp_xcpt_st = T_538;
  assign io_resp_xcpt_if = T_551;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_ptw_req_valid = T_605;
  assign io_ptw_req_bits_addr = r_refill_tag[26:0];
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_store = r_req_store;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign tag_cam_clk = clk;
  assign tag_cam_reset = reset;
  assign tag_cam_io_clear = io_ptw_invalidate;
  assign tag_cam_io_clear_mask = 8'hff;
  assign tag_cam_io_tag = lookup_tag;
  assign tag_cam_io_write = T_169;
  assign tag_cam_io_write_tag = r_refill_tag;
  assign tag_cam_io_write_addr = r_refill_waddr;
  assign tag_ram_T_561_addr = {{2'd0}, 1'h0};
  assign tag_ram_T_561_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_561_data = tag_ram[tag_ram_T_561_addr];
  `else
  assign tag_ram_T_561_data = tag_ram_T_561_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_561_addr];
  `endif
  assign tag_ram_T_563_addr = {{2'd0}, 1'h1};
  assign tag_ram_T_563_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_563_data = tag_ram[tag_ram_T_563_addr];
  `else
  assign tag_ram_T_563_data = tag_ram_T_563_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_563_addr];
  `endif
  assign tag_ram_T_565_addr = {{1'd0}, 2'h2};
  assign tag_ram_T_565_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_565_data = tag_ram[tag_ram_T_565_addr];
  `else
  assign tag_ram_T_565_data = tag_ram_T_565_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_565_addr];
  `endif
  assign tag_ram_T_567_addr = {{1'd0}, 2'h3};
  assign tag_ram_T_567_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_567_data = tag_ram[tag_ram_T_567_addr];
  `else
  assign tag_ram_T_567_data = tag_ram_T_567_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_567_addr];
  `endif
  assign tag_ram_T_569_addr = 3'h4;
  assign tag_ram_T_569_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_569_data = tag_ram[tag_ram_T_569_addr];
  `else
  assign tag_ram_T_569_data = tag_ram_T_569_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_569_addr];
  `endif
  assign tag_ram_T_571_addr = 3'h5;
  assign tag_ram_T_571_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_571_data = tag_ram[tag_ram_T_571_addr];
  `else
  assign tag_ram_T_571_data = tag_ram_T_571_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_571_addr];
  `endif
  assign tag_ram_T_573_addr = 3'h6;
  assign tag_ram_T_573_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_573_data = tag_ram[tag_ram_T_573_addr];
  `else
  assign tag_ram_T_573_data = tag_ram_T_573_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_573_addr];
  `endif
  assign tag_ram_T_575_addr = 3'h7;
  assign tag_ram_T_575_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_575_data = tag_ram[tag_ram_T_575_addr];
  `else
  assign tag_ram_T_575_data = tag_ram_T_575_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_575_addr];
  `endif
  assign tag_ram_T_231_data = io_ptw_resp_bits_pte_ppn;
  assign tag_ram_T_231_addr = r_refill_waddr;
  assign tag_ram_T_231_mask = io_ptw_resp_valid;
  assign tag_ram_T_231_en = io_ptw_resp_valid;
  assign T_167 = io_req_bits_vpn[26:0];
  assign lookup_tag = {io_ptw_ptbr_asid,T_167};
  assign T_168 = state == 2'h2;
  assign T_169 = T_168 & io_ptw_resp_valid;
  assign T_170 = tag_cam_io_hits[7:4];
  assign T_171 = tag_cam_io_hits[3:0];
  assign GEN_145 = {{3'd0}, 1'h0};
  assign T_173 = T_170 != GEN_145;
  assign T_174 = T_170 | T_171;
  assign T_175 = T_174[3:2];
  assign T_176 = T_174[1:0];
  assign GEN_146 = {{1'd0}, 1'h0};
  assign T_178 = T_175 != GEN_146;
  assign T_179 = T_175 | T_176;
  assign T_180 = T_179[1];
  assign T_181 = {T_178,T_180};
  assign tag_hit_addr = {T_173,T_181};
  assign GEN_147 = {{2'd0}, 2'h2};
  assign T_233 = io_ptw_resp_bits_pte_typ >= GEN_147;
  assign T_234 = io_ptw_resp_bits_pte_v & T_233;
  assign T_236 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T_237 = T_234 & T_236;
  assign GEN_0 = T_237;
  assign GEN_148 = {{2'd0}, 1'h0};
  assign GEN_7 = GEN_148 == r_refill_waddr ? GEN_0 : ur_array_0;
  assign GEN_149 = {{2'd0}, 1'h1};
  assign GEN_8 = GEN_149 == r_refill_waddr ? GEN_0 : ur_array_1;
  assign GEN_150 = {{1'd0}, 2'h2};
  assign GEN_9 = GEN_150 == r_refill_waddr ? GEN_0 : ur_array_2;
  assign GEN_151 = {{1'd0}, 2'h3};
  assign GEN_10 = GEN_151 == r_refill_waddr ? GEN_0 : ur_array_3;
  assign GEN_11 = 3'h4 == r_refill_waddr ? GEN_0 : ur_array_4;
  assign GEN_12 = 3'h5 == r_refill_waddr ? GEN_0 : ur_array_5;
  assign GEN_13 = 3'h6 == r_refill_waddr ? GEN_0 : ur_array_6;
  assign GEN_14 = 3'h7 == r_refill_waddr ? GEN_0 : ur_array_7;
  assign T_244 = io_ptw_resp_bits_pte_typ[0];
  assign T_245 = T_237 & T_244;
  assign GEN_1 = T_245;
  assign GEN_15 = GEN_148 == r_refill_waddr ? GEN_1 : uw_array_0;
  assign GEN_16 = GEN_149 == r_refill_waddr ? GEN_1 : uw_array_1;
  assign GEN_17 = GEN_150 == r_refill_waddr ? GEN_1 : uw_array_2;
  assign GEN_18 = GEN_151 == r_refill_waddr ? GEN_1 : uw_array_3;
  assign GEN_19 = 3'h4 == r_refill_waddr ? GEN_1 : uw_array_4;
  assign GEN_20 = 3'h5 == r_refill_waddr ? GEN_1 : uw_array_5;
  assign GEN_21 = 3'h6 == r_refill_waddr ? GEN_1 : uw_array_6;
  assign GEN_22 = 3'h7 == r_refill_waddr ? GEN_1 : uw_array_7;
  assign T_252 = io_ptw_resp_bits_pte_typ[1];
  assign T_253 = T_237 & T_252;
  assign GEN_2 = T_253;
  assign GEN_23 = GEN_148 == r_refill_waddr ? GEN_2 : ux_array_0;
  assign GEN_24 = GEN_149 == r_refill_waddr ? GEN_2 : ux_array_1;
  assign GEN_25 = GEN_150 == r_refill_waddr ? GEN_2 : ux_array_2;
  assign GEN_26 = GEN_151 == r_refill_waddr ? GEN_2 : ux_array_3;
  assign GEN_27 = 3'h4 == r_refill_waddr ? GEN_2 : ux_array_4;
  assign GEN_28 = 3'h5 == r_refill_waddr ? GEN_2 : ux_array_5;
  assign GEN_29 = 3'h6 == r_refill_waddr ? GEN_2 : ux_array_6;
  assign GEN_30 = 3'h7 == r_refill_waddr ? GEN_2 : ux_array_7;
  assign GEN_3 = T_234;
  assign GEN_31 = GEN_148 == r_refill_waddr ? GEN_3 : sr_array_0;
  assign GEN_32 = GEN_149 == r_refill_waddr ? GEN_3 : sr_array_1;
  assign GEN_33 = GEN_150 == r_refill_waddr ? GEN_3 : sr_array_2;
  assign GEN_34 = GEN_151 == r_refill_waddr ? GEN_3 : sr_array_3;
  assign GEN_35 = 3'h4 == r_refill_waddr ? GEN_3 : sr_array_4;
  assign GEN_36 = 3'h5 == r_refill_waddr ? GEN_3 : sr_array_5;
  assign GEN_37 = 3'h6 == r_refill_waddr ? GEN_3 : sr_array_6;
  assign GEN_38 = 3'h7 == r_refill_waddr ? GEN_3 : sr_array_7;
  assign T_261 = T_234 & T_244;
  assign GEN_4 = T_261;
  assign GEN_39 = GEN_148 == r_refill_waddr ? GEN_4 : sw_array_0;
  assign GEN_40 = GEN_149 == r_refill_waddr ? GEN_4 : sw_array_1;
  assign GEN_41 = GEN_150 == r_refill_waddr ? GEN_4 : sw_array_2;
  assign GEN_42 = GEN_151 == r_refill_waddr ? GEN_4 : sw_array_3;
  assign GEN_43 = 3'h4 == r_refill_waddr ? GEN_4 : sw_array_4;
  assign GEN_44 = 3'h5 == r_refill_waddr ? GEN_4 : sw_array_5;
  assign GEN_45 = 3'h6 == r_refill_waddr ? GEN_4 : sw_array_6;
  assign GEN_46 = 3'h7 == r_refill_waddr ? GEN_4 : sw_array_7;
  assign GEN_172 = {{1'd0}, 3'h4};
  assign T_263 = io_ptw_resp_bits_pte_typ >= GEN_172;
  assign T_264 = io_ptw_resp_bits_pte_v & T_263;
  assign T_266 = T_264 & T_252;
  assign GEN_5 = T_266;
  assign GEN_47 = GEN_148 == r_refill_waddr ? GEN_5 : sx_array_0;
  assign GEN_48 = GEN_149 == r_refill_waddr ? GEN_5 : sx_array_1;
  assign GEN_49 = GEN_150 == r_refill_waddr ? GEN_5 : sx_array_2;
  assign GEN_50 = GEN_151 == r_refill_waddr ? GEN_5 : sx_array_3;
  assign GEN_51 = 3'h4 == r_refill_waddr ? GEN_5 : sx_array_4;
  assign GEN_52 = 3'h5 == r_refill_waddr ? GEN_5 : sx_array_5;
  assign GEN_53 = 3'h6 == r_refill_waddr ? GEN_5 : sx_array_6;
  assign GEN_54 = 3'h7 == r_refill_waddr ? GEN_5 : sx_array_7;
  assign GEN_6 = io_ptw_resp_bits_pte_d;
  assign GEN_55 = GEN_148 == r_refill_waddr ? GEN_6 : dirty_array_0;
  assign GEN_56 = GEN_149 == r_refill_waddr ? GEN_6 : dirty_array_1;
  assign GEN_57 = GEN_150 == r_refill_waddr ? GEN_6 : dirty_array_2;
  assign GEN_58 = GEN_151 == r_refill_waddr ? GEN_6 : dirty_array_3;
  assign GEN_59 = 3'h4 == r_refill_waddr ? GEN_6 : dirty_array_4;
  assign GEN_60 = 3'h5 == r_refill_waddr ? GEN_6 : dirty_array_5;
  assign GEN_61 = 3'h6 == r_refill_waddr ? GEN_6 : dirty_array_6;
  assign GEN_62 = 3'h7 == r_refill_waddr ? GEN_6 : dirty_array_7;
  assign GEN_69 = io_ptw_resp_valid ? GEN_7 : ur_array_0;
  assign GEN_70 = io_ptw_resp_valid ? GEN_8 : ur_array_1;
  assign GEN_71 = io_ptw_resp_valid ? GEN_9 : ur_array_2;
  assign GEN_72 = io_ptw_resp_valid ? GEN_10 : ur_array_3;
  assign GEN_73 = io_ptw_resp_valid ? GEN_11 : ur_array_4;
  assign GEN_74 = io_ptw_resp_valid ? GEN_12 : ur_array_5;
  assign GEN_75 = io_ptw_resp_valid ? GEN_13 : ur_array_6;
  assign GEN_76 = io_ptw_resp_valid ? GEN_14 : ur_array_7;
  assign GEN_78 = io_ptw_resp_valid ? GEN_15 : uw_array_0;
  assign GEN_79 = io_ptw_resp_valid ? GEN_16 : uw_array_1;
  assign GEN_80 = io_ptw_resp_valid ? GEN_17 : uw_array_2;
  assign GEN_81 = io_ptw_resp_valid ? GEN_18 : uw_array_3;
  assign GEN_82 = io_ptw_resp_valid ? GEN_19 : uw_array_4;
  assign GEN_83 = io_ptw_resp_valid ? GEN_20 : uw_array_5;
  assign GEN_84 = io_ptw_resp_valid ? GEN_21 : uw_array_6;
  assign GEN_85 = io_ptw_resp_valid ? GEN_22 : uw_array_7;
  assign GEN_87 = io_ptw_resp_valid ? GEN_23 : ux_array_0;
  assign GEN_88 = io_ptw_resp_valid ? GEN_24 : ux_array_1;
  assign GEN_89 = io_ptw_resp_valid ? GEN_25 : ux_array_2;
  assign GEN_90 = io_ptw_resp_valid ? GEN_26 : ux_array_3;
  assign GEN_91 = io_ptw_resp_valid ? GEN_27 : ux_array_4;
  assign GEN_92 = io_ptw_resp_valid ? GEN_28 : ux_array_5;
  assign GEN_93 = io_ptw_resp_valid ? GEN_29 : ux_array_6;
  assign GEN_94 = io_ptw_resp_valid ? GEN_30 : ux_array_7;
  assign GEN_96 = io_ptw_resp_valid ? GEN_31 : sr_array_0;
  assign GEN_97 = io_ptw_resp_valid ? GEN_32 : sr_array_1;
  assign GEN_98 = io_ptw_resp_valid ? GEN_33 : sr_array_2;
  assign GEN_99 = io_ptw_resp_valid ? GEN_34 : sr_array_3;
  assign GEN_100 = io_ptw_resp_valid ? GEN_35 : sr_array_4;
  assign GEN_101 = io_ptw_resp_valid ? GEN_36 : sr_array_5;
  assign GEN_102 = io_ptw_resp_valid ? GEN_37 : sr_array_6;
  assign GEN_103 = io_ptw_resp_valid ? GEN_38 : sr_array_7;
  assign GEN_105 = io_ptw_resp_valid ? GEN_39 : sw_array_0;
  assign GEN_106 = io_ptw_resp_valid ? GEN_40 : sw_array_1;
  assign GEN_107 = io_ptw_resp_valid ? GEN_41 : sw_array_2;
  assign GEN_108 = io_ptw_resp_valid ? GEN_42 : sw_array_3;
  assign GEN_109 = io_ptw_resp_valid ? GEN_43 : sw_array_4;
  assign GEN_110 = io_ptw_resp_valid ? GEN_44 : sw_array_5;
  assign GEN_111 = io_ptw_resp_valid ? GEN_45 : sw_array_6;
  assign GEN_112 = io_ptw_resp_valid ? GEN_46 : sw_array_7;
  assign GEN_114 = io_ptw_resp_valid ? GEN_47 : sx_array_0;
  assign GEN_115 = io_ptw_resp_valid ? GEN_48 : sx_array_1;
  assign GEN_116 = io_ptw_resp_valid ? GEN_49 : sx_array_2;
  assign GEN_117 = io_ptw_resp_valid ? GEN_50 : sx_array_3;
  assign GEN_118 = io_ptw_resp_valid ? GEN_51 : sx_array_4;
  assign GEN_119 = io_ptw_resp_valid ? GEN_52 : sx_array_5;
  assign GEN_120 = io_ptw_resp_valid ? GEN_53 : sx_array_6;
  assign GEN_121 = io_ptw_resp_valid ? GEN_54 : sx_array_7;
  assign GEN_123 = io_ptw_resp_valid ? GEN_55 : dirty_array_0;
  assign GEN_124 = io_ptw_resp_valid ? GEN_56 : dirty_array_1;
  assign GEN_125 = io_ptw_resp_valid ? GEN_57 : dirty_array_2;
  assign GEN_126 = io_ptw_resp_valid ? GEN_58 : dirty_array_3;
  assign GEN_127 = io_ptw_resp_valid ? GEN_59 : dirty_array_4;
  assign GEN_128 = io_ptw_resp_valid ? GEN_60 : dirty_array_5;
  assign GEN_129 = io_ptw_resp_valid ? GEN_61 : dirty_array_6;
  assign GEN_130 = io_ptw_resp_valid ? GEN_62 : dirty_array_7;
  assign T_267 = ~ tag_cam_io_valid_bits;
  assign GEN_181 = {{7'd0}, 1'h0};
  assign T_269 = T_267 == GEN_181;
  assign has_invalid_entry = T_269 == 1'h0;
  assign T_272 = T_267[0];
  assign T_273 = T_267[1];
  assign T_274 = T_267[2];
  assign T_275 = T_267[3];
  assign T_276 = T_267[4];
  assign T_277 = T_267[5];
  assign T_278 = T_267[6];
  assign T_288 = T_278 ? 3'h6 : 3'h7;
  assign T_289 = T_277 ? 3'h5 : T_288;
  assign T_290 = T_276 ? 3'h4 : T_289;
  assign T_291 = T_275 ? {{1'd0}, 2'h3} : T_290;
  assign T_292 = T_274 ? {{1'd0}, 2'h2} : T_291;
  assign T_293 = T_273 ? {{2'd0}, 1'h1} : T_292;
  assign invalid_entry = T_272 ? {{2'd0}, 1'h0} : T_293;
  assign T_297 = T_295 >> 1'h1;
  assign T_298 = T_297[0];
  assign T_299 = {1'h1,T_298};
  assign T_300 = T_295 >> T_299;
  assign T_301 = T_300[0];
  assign T_302 = {T_299,T_301};
  assign T_303 = T_295 >> T_302;
  assign T_304 = T_303[0];
  assign T_305 = {T_302,T_304};
  assign T_306 = T_305[2:0];
  assign repl_waddr = has_invalid_entry ? invalid_entry : T_306;
  assign T_308 = io_req_bits_instruction == 1'h0;
  assign do_mprv = io_ptw_status_mprv & T_308;
  assign priv = do_mprv ? io_ptw_status_mpp : io_ptw_status_prv;
  assign GEN_182 = {{1'd0}, 1'h1};
  assign priv_s = priv == GEN_182;
  assign T_311 = priv <= GEN_182;
  assign T_313 = io_ptw_status_debug == 1'h0;
  assign priv_uses_vm = T_311 & T_313;
  assign T_320 = {ur_array_1,ur_array_0};
  assign T_321 = {ur_array_3,ur_array_2};
  assign T_322 = {T_321,T_320};
  assign T_323 = {ur_array_5,ur_array_4};
  assign T_324 = {ur_array_7,ur_array_6};
  assign T_325 = {T_324,T_323};
  assign ur_bits = {T_325,T_322};
  assign T_327 = io_ptw_status_pum ? ur_bits : {{7'd0}, 1'h0};
  assign pum_ok = ~ T_327;
  assign T_328 = {sr_array_1,sr_array_0};
  assign T_329 = {sr_array_3,sr_array_2};
  assign T_330 = {T_329,T_328};
  assign T_331 = {sr_array_5,sr_array_4};
  assign T_332 = {sr_array_7,sr_array_6};
  assign T_333 = {T_332,T_331};
  assign T_334 = {T_333,T_330};
  assign T_335 = T_334 & pum_ok;
  assign r_array = priv_s ? T_335 : ur_bits;
  assign T_336 = {sw_array_1,sw_array_0};
  assign T_337 = {sw_array_3,sw_array_2};
  assign T_338 = {T_337,T_336};
  assign T_339 = {sw_array_5,sw_array_4};
  assign T_340 = {sw_array_7,sw_array_6};
  assign T_341 = {T_340,T_339};
  assign T_342 = {T_341,T_338};
  assign T_343 = T_342 & pum_ok;
  assign T_344 = {uw_array_1,uw_array_0};
  assign T_345 = {uw_array_3,uw_array_2};
  assign T_346 = {T_345,T_344};
  assign T_347 = {uw_array_5,uw_array_4};
  assign T_348 = {uw_array_7,uw_array_6};
  assign T_349 = {T_348,T_347};
  assign T_350 = {T_349,T_346};
  assign w_array = priv_s ? T_343 : T_350;
  assign T_351 = {sx_array_1,sx_array_0};
  assign T_352 = {sx_array_3,sx_array_2};
  assign T_353 = {T_352,T_351};
  assign T_354 = {sx_array_5,sx_array_4};
  assign T_355 = {sx_array_7,sx_array_6};
  assign T_356 = {T_355,T_354};
  assign T_357 = {T_356,T_353};
  assign T_358 = {ux_array_1,ux_array_0};
  assign T_359 = {ux_array_3,ux_array_2};
  assign T_360 = {T_359,T_358};
  assign T_361 = {ux_array_5,ux_array_4};
  assign T_362 = {ux_array_7,ux_array_6};
  assign T_363 = {T_362,T_361};
  assign T_364 = {T_363,T_360};
  assign x_array = priv_s ? T_357 : T_364;
  assign T_366 = io_ptw_status_vm[3];
  assign T_368 = T_366 & priv_uses_vm;
  assign T_370 = io_req_bits_passthrough == 1'h0;
  assign vm_enabled = T_368 & T_370;
  assign T_371 = io_req_bits_vpn[27];
  assign T_372 = io_req_bits_vpn[26];
  assign bad_va = T_371 != T_372;
  assign T_373 = {dirty_array_1,dirty_array_0};
  assign T_374 = {dirty_array_3,dirty_array_2};
  assign T_375 = {T_374,T_373};
  assign T_376 = {dirty_array_5,dirty_array_4};
  assign T_377 = {dirty_array_7,dirty_array_6};
  assign T_378 = {T_377,T_376};
  assign T_379 = {T_378,T_375};
  assign T_381 = io_req_bits_store ? w_array : {{7'd0}, 1'h0};
  assign T_382 = ~ T_381;
  assign T_383 = T_379 | T_382;
  assign tag_hits = tag_cam_io_hits & T_383;
  assign tag_hit = tag_hits != GEN_181;
  assign tlb_hit = vm_enabled & tag_hit;
  assign T_386 = tag_hit == 1'h0;
  assign T_387 = vm_enabled & T_386;
  assign T_389 = bad_va == 1'h0;
  assign tlb_miss = T_387 & T_389;
  assign T_390 = io_req_valid & tlb_hit;
  assign T_405 = tag_hit_addr[2];
  assign GEN_187 = {{1'd0}, 8'h1};
  assign T_407 = GEN_187 << 1'h1;
  assign T_408 = T_407[7:0];
  assign T_409 = ~ T_408;
  assign T_410 = T_295 & T_409;
  assign T_412 = T_405 ? {{7'd0}, 1'h0} : T_408;
  assign T_413 = T_410 | T_412;
  assign T_414 = {1'h1,T_405};
  assign T_415 = tag_hit_addr[1];
  assign GEN_188 = {{3'd0}, 8'h1};
  assign T_417 = GEN_188 << T_414;
  assign T_418 = T_417[7:0];
  assign T_419 = ~ T_418;
  assign T_420 = T_413 & T_419;
  assign T_422 = T_415 ? {{7'd0}, 1'h0} : T_418;
  assign T_423 = T_420 | T_422;
  assign T_424 = {T_414,T_415};
  assign T_425 = tag_hit_addr[0];
  assign GEN_189 = {{7'd0}, 8'h1};
  assign T_427 = GEN_189 << T_424;
  assign T_428 = T_427[7:0];
  assign T_429 = ~ T_428;
  assign T_430 = T_423 & T_429;
  assign T_432 = T_425 ? {{7'd0}, 1'h0} : T_428;
  assign T_433 = T_430 | T_432;
  assign GEN_131 = T_390 ? T_433 : T_295;
  assign paddr = {io_resp_ppn,12'h0};
  assign GEN_190 = {{19'd0}, 13'h1000};
  assign T_439 = paddr < GEN_190;
  assign T_443 = T_439 ? 3'h7 : {{2'd0}, 1'h0};
  assign T_445 = GEN_190 <= paddr;
  assign GEN_192 = {{18'd0}, 14'h2000};
  assign T_447 = paddr < GEN_192;
  assign T_448 = T_445 & T_447;
  assign T_451 = T_448 ? 3'h5 : {{2'd0}, 1'h0};
  assign T_453 = GEN_192 <= paddr;
  assign GEN_194 = {{17'd0}, 15'h4000};
  assign T_455 = paddr < GEN_194;
  assign T_456 = T_453 & T_455;
  assign T_459 = T_456 ? 3'h7 : {{2'd0}, 1'h0};
  assign GEN_195 = {{1'd0}, 31'h40000000};
  assign T_461 = GEN_195 <= paddr;
  assign GEN_196 = {{1'd0}, 31'h44000000};
  assign T_463 = paddr < GEN_196;
  assign T_464 = T_461 & T_463;
  assign T_467 = T_464 ? 3'h3 : {{2'd0}, 1'h0};
  assign T_469 = GEN_196 <= paddr;
  assign GEN_198 = {{1'd0}, 31'h48000000};
  assign T_471 = paddr < GEN_198;
  assign T_472 = T_469 & T_471;
  assign T_475 = T_472 ? 3'h3 : {{2'd0}, 1'h0};
  assign GEN_199 = {{1'd0}, 31'h60000000};
  assign T_477 = GEN_199 <= paddr;
  assign T_479 = paddr < 32'h80000000;
  assign T_480 = T_477 & T_479;
  assign T_483 = T_480 ? 3'h7 : {{2'd0}, 1'h0};
  assign T_485 = 32'h80000000 <= paddr;
  assign T_491 = T_485 ? 3'h7 : {{2'd0}, 1'h0};
  assign T_496 = T_443 | T_451;
  assign T_497 = T_496 | T_459;
  assign T_498 = T_497 | T_467;
  assign T_499 = T_498 | T_475;
  assign T_500 = T_499 | T_483;
  assign T_501 = T_500 | T_491;
  assign addr_prot_x = T_511;
  assign addr_prot_w = T_510;
  assign addr_prot_r = T_509;
  assign T_509 = T_501[0];
  assign T_510 = T_501[1];
  assign T_511 = T_501[2];
  assign T_512 = state == 2'h0;
  assign T_514 = tlb_miss == 1'h0;
  assign T_516 = addr_prot_r == 1'h0;
  assign T_517 = T_514 & T_516;
  assign T_518 = bad_va | T_517;
  assign T_519 = r_array & tag_cam_io_hits;
  assign T_521 = T_519 != GEN_181;
  assign T_523 = T_521 == 1'h0;
  assign T_524 = tlb_hit & T_523;
  assign T_525 = T_518 | T_524;
  assign T_529 = addr_prot_w == 1'h0;
  assign T_530 = T_514 & T_529;
  assign T_531 = bad_va | T_530;
  assign T_532 = w_array & tag_cam_io_hits;
  assign T_534 = T_532 != GEN_181;
  assign T_536 = T_534 == 1'h0;
  assign T_537 = tlb_hit & T_536;
  assign T_538 = T_531 | T_537;
  assign T_542 = addr_prot_x == 1'h0;
  assign T_543 = T_514 & T_542;
  assign T_544 = bad_va | T_543;
  assign T_545 = x_array & tag_cam_io_hits;
  assign T_547 = T_545 != GEN_181;
  assign T_549 = T_547 == 1'h0;
  assign T_550 = tlb_hit & T_549;
  assign T_551 = T_544 | T_550;
  assign T_552 = tag_cam_io_hits[0];
  assign T_553 = tag_cam_io_hits[1];
  assign T_554 = tag_cam_io_hits[2];
  assign T_555 = tag_cam_io_hits[3];
  assign T_556 = tag_cam_io_hits[4];
  assign T_557 = tag_cam_io_hits[5];
  assign T_558 = tag_cam_io_hits[6];
  assign T_559 = tag_cam_io_hits[7];
  assign T_577 = T_552 ? tag_ram_T_561_data : {{19'd0}, 1'h0};
  assign T_579 = T_553 ? tag_ram_T_563_data : {{19'd0}, 1'h0};
  assign T_581 = T_554 ? tag_ram_T_565_data : {{19'd0}, 1'h0};
  assign T_583 = T_555 ? tag_ram_T_567_data : {{19'd0}, 1'h0};
  assign T_585 = T_556 ? tag_ram_T_569_data : {{19'd0}, 1'h0};
  assign T_587 = T_557 ? tag_ram_T_571_data : {{19'd0}, 1'h0};
  assign T_589 = T_558 ? tag_ram_T_573_data : {{19'd0}, 1'h0};
  assign T_591 = T_559 ? tag_ram_T_575_data : {{19'd0}, 1'h0};
  assign T_593 = T_577 | T_579;
  assign T_594 = T_593 | T_581;
  assign T_595 = T_594 | T_583;
  assign T_596 = T_595 | T_585;
  assign T_597 = T_596 | T_587;
  assign T_598 = T_597 | T_589;
  assign T_599 = T_598 | T_591;
  assign T_600 = T_599;
  assign T_601 = io_req_bits_vpn[19:0];
  assign T_602 = vm_enabled ? T_600 : T_601;
  assign T_605 = state == 2'h1;
  assign T_606 = io_req_ready & io_req_valid;
  assign T_607 = T_606 & tlb_miss;
  assign GEN_132 = T_607 ? 2'h1 : state;
  assign GEN_133 = T_607 ? lookup_tag : r_refill_tag;
  assign GEN_134 = T_607 ? repl_waddr : r_refill_waddr;
  assign GEN_135 = T_607 ? io_req_bits_vpn : r_req_vpn;
  assign GEN_136 = T_607 ? io_req_bits_passthrough : r_req_passthrough;
  assign GEN_137 = T_607 ? io_req_bits_instruction : r_req_instruction;
  assign GEN_138 = T_607 ? io_req_bits_store : r_req_store;
  assign GEN_139 = io_ptw_invalidate ? 2'h0 : GEN_132;
  assign GEN_140 = io_ptw_invalidate ? 2'h3 : 2'h2;
  assign GEN_141 = io_ptw_req_ready ? GEN_140 : GEN_139;
  assign GEN_142 = T_605 ? GEN_141 : GEN_132;
  assign T_610 = T_168 & io_ptw_invalidate;
  assign GEN_143 = T_610 ? 2'h3 : GEN_142;
  assign GEN_144 = io_ptw_resp_valid ? 2'h0 : GEN_143;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_63 = {1{$random}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    tag_ram[initvar] = GEN_63[19:0];
  GEN_64 = {1{$random}};
  state = GEN_64[1:0];
  GEN_65 = {2{$random}};
  r_refill_tag = GEN_65[33:0];
  GEN_66 = {1{$random}};
  r_refill_waddr = GEN_66[2:0];
  GEN_67 = {1{$random}};
  r_req_vpn = GEN_67[27:0];
  GEN_68 = {1{$random}};
  r_req_passthrough = GEN_68[0:0];
  GEN_77 = {1{$random}};
  r_req_instruction = GEN_77[0:0];
  GEN_86 = {1{$random}};
  r_req_store = GEN_86[0:0];
  GEN_95 = {1{$random}};
  ur_array_0 = GEN_95[0:0];
  GEN_104 = {1{$random}};
  ur_array_1 = GEN_104[0:0];
  GEN_113 = {1{$random}};
  ur_array_2 = GEN_113[0:0];
  GEN_122 = {1{$random}};
  ur_array_3 = GEN_122[0:0];
  GEN_152 = {1{$random}};
  ur_array_4 = GEN_152[0:0];
  GEN_153 = {1{$random}};
  ur_array_5 = GEN_153[0:0];
  GEN_154 = {1{$random}};
  ur_array_6 = GEN_154[0:0];
  GEN_155 = {1{$random}};
  ur_array_7 = GEN_155[0:0];
  GEN_156 = {1{$random}};
  uw_array_0 = GEN_156[0:0];
  GEN_157 = {1{$random}};
  uw_array_1 = GEN_157[0:0];
  GEN_158 = {1{$random}};
  uw_array_2 = GEN_158[0:0];
  GEN_159 = {1{$random}};
  uw_array_3 = GEN_159[0:0];
  GEN_160 = {1{$random}};
  uw_array_4 = GEN_160[0:0];
  GEN_161 = {1{$random}};
  uw_array_5 = GEN_161[0:0];
  GEN_162 = {1{$random}};
  uw_array_6 = GEN_162[0:0];
  GEN_163 = {1{$random}};
  uw_array_7 = GEN_163[0:0];
  GEN_164 = {1{$random}};
  ux_array_0 = GEN_164[0:0];
  GEN_165 = {1{$random}};
  ux_array_1 = GEN_165[0:0];
  GEN_166 = {1{$random}};
  ux_array_2 = GEN_166[0:0];
  GEN_167 = {1{$random}};
  ux_array_3 = GEN_167[0:0];
  GEN_168 = {1{$random}};
  ux_array_4 = GEN_168[0:0];
  GEN_169 = {1{$random}};
  ux_array_5 = GEN_169[0:0];
  GEN_170 = {1{$random}};
  ux_array_6 = GEN_170[0:0];
  GEN_171 = {1{$random}};
  ux_array_7 = GEN_171[0:0];
  GEN_173 = {1{$random}};
  sr_array_0 = GEN_173[0:0];
  GEN_174 = {1{$random}};
  sr_array_1 = GEN_174[0:0];
  GEN_175 = {1{$random}};
  sr_array_2 = GEN_175[0:0];
  GEN_176 = {1{$random}};
  sr_array_3 = GEN_176[0:0];
  GEN_177 = {1{$random}};
  sr_array_4 = GEN_177[0:0];
  GEN_178 = {1{$random}};
  sr_array_5 = GEN_178[0:0];
  GEN_179 = {1{$random}};
  sr_array_6 = GEN_179[0:0];
  GEN_180 = {1{$random}};
  sr_array_7 = GEN_180[0:0];
  GEN_183 = {1{$random}};
  sw_array_0 = GEN_183[0:0];
  GEN_184 = {1{$random}};
  sw_array_1 = GEN_184[0:0];
  GEN_185 = {1{$random}};
  sw_array_2 = GEN_185[0:0];
  GEN_186 = {1{$random}};
  sw_array_3 = GEN_186[0:0];
  GEN_191 = {1{$random}};
  sw_array_4 = GEN_191[0:0];
  GEN_193 = {1{$random}};
  sw_array_5 = GEN_193[0:0];
  GEN_197 = {1{$random}};
  sw_array_6 = GEN_197[0:0];
  GEN_200 = {1{$random}};
  sw_array_7 = GEN_200[0:0];
  GEN_201 = {1{$random}};
  sx_array_0 = GEN_201[0:0];
  GEN_202 = {1{$random}};
  sx_array_1 = GEN_202[0:0];
  GEN_203 = {1{$random}};
  sx_array_2 = GEN_203[0:0];
  GEN_204 = {1{$random}};
  sx_array_3 = GEN_204[0:0];
  GEN_205 = {1{$random}};
  sx_array_4 = GEN_205[0:0];
  GEN_206 = {1{$random}};
  sx_array_5 = GEN_206[0:0];
  GEN_207 = {1{$random}};
  sx_array_6 = GEN_207[0:0];
  GEN_208 = {1{$random}};
  sx_array_7 = GEN_208[0:0];
  GEN_209 = {1{$random}};
  dirty_array_0 = GEN_209[0:0];
  GEN_210 = {1{$random}};
  dirty_array_1 = GEN_210[0:0];
  GEN_211 = {1{$random}};
  dirty_array_2 = GEN_211[0:0];
  GEN_212 = {1{$random}};
  dirty_array_3 = GEN_212[0:0];
  GEN_213 = {1{$random}};
  dirty_array_4 = GEN_213[0:0];
  GEN_214 = {1{$random}};
  dirty_array_5 = GEN_214[0:0];
  GEN_215 = {1{$random}};
  dirty_array_6 = GEN_215[0:0];
  GEN_216 = {1{$random}};
  dirty_array_7 = GEN_216[0:0];
  GEN_217 = {1{$random}};
  T_295 = GEN_217[7:0];
  end
`endif
  always @(posedge clk) begin
    if(tag_ram_T_231_en & tag_ram_T_231_mask) begin
      tag_ram[tag_ram_T_231_addr] <= tag_ram_T_231_data;
    end
    if(reset) begin
      state <= 2'h0;
    end else begin
      if(io_ptw_resp_valid) begin
        state <= 2'h0;
      end else begin
        if(T_610) begin
          state <= 2'h3;
        end else begin
          if(T_605) begin
            if(io_ptw_req_ready) begin
              if(io_ptw_invalidate) begin
                state <= 2'h3;
              end else begin
                state <= 2'h2;
              end
            end else begin
              if(io_ptw_invalidate) begin
                state <= 2'h0;
              end else begin
                if(T_607) begin
                  state <= 2'h1;
                end
              end
            end
          end else begin
            if(T_607) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_607) begin
        r_refill_tag <= lookup_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_607) begin
        if(has_invalid_entry) begin
          if(T_272) begin
            r_refill_waddr <= {{2'd0}, 1'h0};
          end else begin
            if(T_273) begin
              r_refill_waddr <= {{2'd0}, 1'h1};
            end else begin
              if(T_274) begin
                r_refill_waddr <= {{1'd0}, 2'h2};
              end else begin
                if(T_275) begin
                  r_refill_waddr <= {{1'd0}, 2'h3};
                end else begin
                  if(T_276) begin
                    r_refill_waddr <= 3'h4;
                  end else begin
                    if(T_277) begin
                      r_refill_waddr <= 3'h5;
                    end else begin
                      if(T_278) begin
                        r_refill_waddr <= 3'h6;
                      end else begin
                        r_refill_waddr <= 3'h7;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          r_refill_waddr <= T_306;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_607) begin
        r_req_vpn <= io_req_bits_vpn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_607) begin
        r_req_passthrough <= io_req_bits_passthrough;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_607) begin
        r_req_instruction <= io_req_bits_instruction;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_607) begin
        r_req_store <= io_req_bits_store;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_148 == r_refill_waddr) begin
          ur_array_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_149 == r_refill_waddr) begin
          ur_array_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_150 == r_refill_waddr) begin
          ur_array_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_151 == r_refill_waddr) begin
          ur_array_3 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          ur_array_4 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          ur_array_5 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          ur_array_6 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          ur_array_7 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_148 == r_refill_waddr) begin
          uw_array_0 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_149 == r_refill_waddr) begin
          uw_array_1 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_150 == r_refill_waddr) begin
          uw_array_2 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_151 == r_refill_waddr) begin
          uw_array_3 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          uw_array_4 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          uw_array_5 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          uw_array_6 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          uw_array_7 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_148 == r_refill_waddr) begin
          ux_array_0 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_149 == r_refill_waddr) begin
          ux_array_1 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_150 == r_refill_waddr) begin
          ux_array_2 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_151 == r_refill_waddr) begin
          ux_array_3 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          ux_array_4 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          ux_array_5 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          ux_array_6 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          ux_array_7 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_148 == r_refill_waddr) begin
          sr_array_0 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_149 == r_refill_waddr) begin
          sr_array_1 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_150 == r_refill_waddr) begin
          sr_array_2 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_151 == r_refill_waddr) begin
          sr_array_3 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          sr_array_4 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          sr_array_5 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          sr_array_6 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          sr_array_7 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_148 == r_refill_waddr) begin
          sw_array_0 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_149 == r_refill_waddr) begin
          sw_array_1 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_150 == r_refill_waddr) begin
          sw_array_2 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_151 == r_refill_waddr) begin
          sw_array_3 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          sw_array_4 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          sw_array_5 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          sw_array_6 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          sw_array_7 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_148 == r_refill_waddr) begin
          sx_array_0 <= GEN_5;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_149 == r_refill_waddr) begin
          sx_array_1 <= GEN_5;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_150 == r_refill_waddr) begin
          sx_array_2 <= GEN_5;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_151 == r_refill_waddr) begin
          sx_array_3 <= GEN_5;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          sx_array_4 <= GEN_5;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          sx_array_5 <= GEN_5;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          sx_array_6 <= GEN_5;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          sx_array_7 <= GEN_5;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_148 == r_refill_waddr) begin
          dirty_array_0 <= GEN_6;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_149 == r_refill_waddr) begin
          dirty_array_1 <= GEN_6;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_150 == r_refill_waddr) begin
          dirty_array_2 <= GEN_6;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(GEN_151 == r_refill_waddr) begin
          dirty_array_3 <= GEN_6;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          dirty_array_4 <= GEN_6;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          dirty_array_5 <= GEN_6;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          dirty_array_6 <= GEN_6;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          dirty_array_7 <= GEN_6;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_390) begin
        T_295 <= T_433;
      end
    end
  end
endmodule
module BTB(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [38:0] io_req_bits_addr,
  output  io_resp_valid,
  output  io_resp_bits_taken,
  output  io_resp_bits_mask,
  output  io_resp_bits_bridx,
  output [38:0] io_resp_bits_target,
  output [5:0] io_resp_bits_entry,
  output [6:0] io_resp_bits_bht_history,
  output [1:0] io_resp_bits_bht_value,
  input   io_btb_update_valid,
  input   io_btb_update_bits_prediction_valid,
  input   io_btb_update_bits_prediction_bits_taken,
  input   io_btb_update_bits_prediction_bits_mask,
  input   io_btb_update_bits_prediction_bits_bridx,
  input  [38:0] io_btb_update_bits_prediction_bits_target,
  input  [5:0] io_btb_update_bits_prediction_bits_entry,
  input  [6:0] io_btb_update_bits_prediction_bits_bht_history,
  input  [1:0] io_btb_update_bits_prediction_bits_bht_value,
  input  [38:0] io_btb_update_bits_pc,
  input  [38:0] io_btb_update_bits_target,
  input   io_btb_update_bits_taken,
  input   io_btb_update_bits_isJump,
  input   io_btb_update_bits_isReturn,
  input  [38:0] io_btb_update_bits_br_pc,
  input   io_bht_update_valid,
  input   io_bht_update_bits_prediction_valid,
  input   io_bht_update_bits_prediction_bits_taken,
  input   io_bht_update_bits_prediction_bits_mask,
  input   io_bht_update_bits_prediction_bits_bridx,
  input  [38:0] io_bht_update_bits_prediction_bits_target,
  input  [5:0] io_bht_update_bits_prediction_bits_entry,
  input  [6:0] io_bht_update_bits_prediction_bits_bht_history,
  input  [1:0] io_bht_update_bits_prediction_bits_bht_value,
  input  [38:0] io_bht_update_bits_pc,
  input   io_bht_update_bits_taken,
  input   io_bht_update_bits_mispredict,
  input   io_ras_update_valid,
  input   io_ras_update_bits_isCall,
  input   io_ras_update_bits_isReturn,
  input  [38:0] io_ras_update_bits_returnAddr,
  input   io_ras_update_bits_prediction_valid,
  input   io_ras_update_bits_prediction_bits_taken,
  input   io_ras_update_bits_prediction_bits_mask,
  input   io_ras_update_bits_prediction_bits_bridx,
  input  [38:0] io_ras_update_bits_prediction_bits_target,
  input  [5:0] io_ras_update_bits_prediction_bits_entry,
  input  [6:0] io_ras_update_bits_prediction_bits_bht_history,
  input  [1:0] io_ras_update_bits_prediction_bits_bht_value,
  input   io_invalidate
);
  reg [61:0] idxValid;
  reg [63:0] GEN_146;
  reg [11:0] idxs [0:61];
  reg [31:0] GEN_147;
  wire [11:0] idxs_T_1431_data;
  wire [5:0] idxs_T_1431_addr;
  wire  idxs_T_1431_en;
  wire [11:0] idxs_T_1434_data;
  wire [5:0] idxs_T_1434_addr;
  wire  idxs_T_1434_en;
  wire [11:0] idxs_T_1437_data;
  wire [5:0] idxs_T_1437_addr;
  wire  idxs_T_1437_en;
  wire [11:0] idxs_T_1440_data;
  wire [5:0] idxs_T_1440_addr;
  wire  idxs_T_1440_en;
  wire [11:0] idxs_T_1443_data;
  wire [5:0] idxs_T_1443_addr;
  wire  idxs_T_1443_en;
  wire [11:0] idxs_T_1446_data;
  wire [5:0] idxs_T_1446_addr;
  wire  idxs_T_1446_en;
  wire [11:0] idxs_T_1449_data;
  wire [5:0] idxs_T_1449_addr;
  wire  idxs_T_1449_en;
  wire [11:0] idxs_T_1452_data;
  wire [5:0] idxs_T_1452_addr;
  wire  idxs_T_1452_en;
  wire [11:0] idxs_T_1455_data;
  wire [5:0] idxs_T_1455_addr;
  wire  idxs_T_1455_en;
  wire [11:0] idxs_T_1458_data;
  wire [5:0] idxs_T_1458_addr;
  wire  idxs_T_1458_en;
  wire [11:0] idxs_T_1461_data;
  wire [5:0] idxs_T_1461_addr;
  wire  idxs_T_1461_en;
  wire [11:0] idxs_T_1464_data;
  wire [5:0] idxs_T_1464_addr;
  wire  idxs_T_1464_en;
  wire [11:0] idxs_T_1467_data;
  wire [5:0] idxs_T_1467_addr;
  wire  idxs_T_1467_en;
  wire [11:0] idxs_T_1470_data;
  wire [5:0] idxs_T_1470_addr;
  wire  idxs_T_1470_en;
  wire [11:0] idxs_T_1473_data;
  wire [5:0] idxs_T_1473_addr;
  wire  idxs_T_1473_en;
  wire [11:0] idxs_T_1476_data;
  wire [5:0] idxs_T_1476_addr;
  wire  idxs_T_1476_en;
  wire [11:0] idxs_T_1479_data;
  wire [5:0] idxs_T_1479_addr;
  wire  idxs_T_1479_en;
  wire [11:0] idxs_T_1482_data;
  wire [5:0] idxs_T_1482_addr;
  wire  idxs_T_1482_en;
  wire [11:0] idxs_T_1485_data;
  wire [5:0] idxs_T_1485_addr;
  wire  idxs_T_1485_en;
  wire [11:0] idxs_T_1488_data;
  wire [5:0] idxs_T_1488_addr;
  wire  idxs_T_1488_en;
  wire [11:0] idxs_T_1491_data;
  wire [5:0] idxs_T_1491_addr;
  wire  idxs_T_1491_en;
  wire [11:0] idxs_T_1494_data;
  wire [5:0] idxs_T_1494_addr;
  wire  idxs_T_1494_en;
  wire [11:0] idxs_T_1497_data;
  wire [5:0] idxs_T_1497_addr;
  wire  idxs_T_1497_en;
  wire [11:0] idxs_T_1500_data;
  wire [5:0] idxs_T_1500_addr;
  wire  idxs_T_1500_en;
  wire [11:0] idxs_T_1503_data;
  wire [5:0] idxs_T_1503_addr;
  wire  idxs_T_1503_en;
  wire [11:0] idxs_T_1506_data;
  wire [5:0] idxs_T_1506_addr;
  wire  idxs_T_1506_en;
  wire [11:0] idxs_T_1509_data;
  wire [5:0] idxs_T_1509_addr;
  wire  idxs_T_1509_en;
  wire [11:0] idxs_T_1512_data;
  wire [5:0] idxs_T_1512_addr;
  wire  idxs_T_1512_en;
  wire [11:0] idxs_T_1515_data;
  wire [5:0] idxs_T_1515_addr;
  wire  idxs_T_1515_en;
  wire [11:0] idxs_T_1518_data;
  wire [5:0] idxs_T_1518_addr;
  wire  idxs_T_1518_en;
  wire [11:0] idxs_T_1521_data;
  wire [5:0] idxs_T_1521_addr;
  wire  idxs_T_1521_en;
  wire [11:0] idxs_T_1524_data;
  wire [5:0] idxs_T_1524_addr;
  wire  idxs_T_1524_en;
  wire [11:0] idxs_T_1527_data;
  wire [5:0] idxs_T_1527_addr;
  wire  idxs_T_1527_en;
  wire [11:0] idxs_T_1530_data;
  wire [5:0] idxs_T_1530_addr;
  wire  idxs_T_1530_en;
  wire [11:0] idxs_T_1533_data;
  wire [5:0] idxs_T_1533_addr;
  wire  idxs_T_1533_en;
  wire [11:0] idxs_T_1536_data;
  wire [5:0] idxs_T_1536_addr;
  wire  idxs_T_1536_en;
  wire [11:0] idxs_T_1539_data;
  wire [5:0] idxs_T_1539_addr;
  wire  idxs_T_1539_en;
  wire [11:0] idxs_T_1542_data;
  wire [5:0] idxs_T_1542_addr;
  wire  idxs_T_1542_en;
  wire [11:0] idxs_T_1545_data;
  wire [5:0] idxs_T_1545_addr;
  wire  idxs_T_1545_en;
  wire [11:0] idxs_T_1548_data;
  wire [5:0] idxs_T_1548_addr;
  wire  idxs_T_1548_en;
  wire [11:0] idxs_T_1551_data;
  wire [5:0] idxs_T_1551_addr;
  wire  idxs_T_1551_en;
  wire [11:0] idxs_T_1554_data;
  wire [5:0] idxs_T_1554_addr;
  wire  idxs_T_1554_en;
  wire [11:0] idxs_T_1557_data;
  wire [5:0] idxs_T_1557_addr;
  wire  idxs_T_1557_en;
  wire [11:0] idxs_T_1560_data;
  wire [5:0] idxs_T_1560_addr;
  wire  idxs_T_1560_en;
  wire [11:0] idxs_T_1563_data;
  wire [5:0] idxs_T_1563_addr;
  wire  idxs_T_1563_en;
  wire [11:0] idxs_T_1566_data;
  wire [5:0] idxs_T_1566_addr;
  wire  idxs_T_1566_en;
  wire [11:0] idxs_T_1569_data;
  wire [5:0] idxs_T_1569_addr;
  wire  idxs_T_1569_en;
  wire [11:0] idxs_T_1572_data;
  wire [5:0] idxs_T_1572_addr;
  wire  idxs_T_1572_en;
  wire [11:0] idxs_T_1575_data;
  wire [5:0] idxs_T_1575_addr;
  wire  idxs_T_1575_en;
  wire [11:0] idxs_T_1578_data;
  wire [5:0] idxs_T_1578_addr;
  wire  idxs_T_1578_en;
  wire [11:0] idxs_T_1581_data;
  wire [5:0] idxs_T_1581_addr;
  wire  idxs_T_1581_en;
  wire [11:0] idxs_T_1584_data;
  wire [5:0] idxs_T_1584_addr;
  wire  idxs_T_1584_en;
  wire [11:0] idxs_T_1587_data;
  wire [5:0] idxs_T_1587_addr;
  wire  idxs_T_1587_en;
  wire [11:0] idxs_T_1590_data;
  wire [5:0] idxs_T_1590_addr;
  wire  idxs_T_1590_en;
  wire [11:0] idxs_T_1593_data;
  wire [5:0] idxs_T_1593_addr;
  wire  idxs_T_1593_en;
  wire [11:0] idxs_T_1596_data;
  wire [5:0] idxs_T_1596_addr;
  wire  idxs_T_1596_en;
  wire [11:0] idxs_T_1599_data;
  wire [5:0] idxs_T_1599_addr;
  wire  idxs_T_1599_en;
  wire [11:0] idxs_T_1602_data;
  wire [5:0] idxs_T_1602_addr;
  wire  idxs_T_1602_en;
  wire [11:0] idxs_T_1605_data;
  wire [5:0] idxs_T_1605_addr;
  wire  idxs_T_1605_en;
  wire [11:0] idxs_T_1608_data;
  wire [5:0] idxs_T_1608_addr;
  wire  idxs_T_1608_en;
  wire [11:0] idxs_T_1611_data;
  wire [5:0] idxs_T_1611_addr;
  wire  idxs_T_1611_en;
  wire [11:0] idxs_T_1614_data;
  wire [5:0] idxs_T_1614_addr;
  wire  idxs_T_1614_en;
  wire [11:0] idxs_T_1972_data;
  wire [5:0] idxs_T_1972_addr;
  wire  idxs_T_1972_en;
  wire [11:0] idxs_T_1975_data;
  wire [5:0] idxs_T_1975_addr;
  wire  idxs_T_1975_en;
  wire [11:0] idxs_T_1978_data;
  wire [5:0] idxs_T_1978_addr;
  wire  idxs_T_1978_en;
  wire [11:0] idxs_T_1981_data;
  wire [5:0] idxs_T_1981_addr;
  wire  idxs_T_1981_en;
  wire [11:0] idxs_T_1984_data;
  wire [5:0] idxs_T_1984_addr;
  wire  idxs_T_1984_en;
  wire [11:0] idxs_T_1987_data;
  wire [5:0] idxs_T_1987_addr;
  wire  idxs_T_1987_en;
  wire [11:0] idxs_T_1990_data;
  wire [5:0] idxs_T_1990_addr;
  wire  idxs_T_1990_en;
  wire [11:0] idxs_T_1993_data;
  wire [5:0] idxs_T_1993_addr;
  wire  idxs_T_1993_en;
  wire [11:0] idxs_T_1996_data;
  wire [5:0] idxs_T_1996_addr;
  wire  idxs_T_1996_en;
  wire [11:0] idxs_T_1999_data;
  wire [5:0] idxs_T_1999_addr;
  wire  idxs_T_1999_en;
  wire [11:0] idxs_T_2002_data;
  wire [5:0] idxs_T_2002_addr;
  wire  idxs_T_2002_en;
  wire [11:0] idxs_T_2005_data;
  wire [5:0] idxs_T_2005_addr;
  wire  idxs_T_2005_en;
  wire [11:0] idxs_T_2008_data;
  wire [5:0] idxs_T_2008_addr;
  wire  idxs_T_2008_en;
  wire [11:0] idxs_T_2011_data;
  wire [5:0] idxs_T_2011_addr;
  wire  idxs_T_2011_en;
  wire [11:0] idxs_T_2014_data;
  wire [5:0] idxs_T_2014_addr;
  wire  idxs_T_2014_en;
  wire [11:0] idxs_T_2017_data;
  wire [5:0] idxs_T_2017_addr;
  wire  idxs_T_2017_en;
  wire [11:0] idxs_T_2020_data;
  wire [5:0] idxs_T_2020_addr;
  wire  idxs_T_2020_en;
  wire [11:0] idxs_T_2023_data;
  wire [5:0] idxs_T_2023_addr;
  wire  idxs_T_2023_en;
  wire [11:0] idxs_T_2026_data;
  wire [5:0] idxs_T_2026_addr;
  wire  idxs_T_2026_en;
  wire [11:0] idxs_T_2029_data;
  wire [5:0] idxs_T_2029_addr;
  wire  idxs_T_2029_en;
  wire [11:0] idxs_T_2032_data;
  wire [5:0] idxs_T_2032_addr;
  wire  idxs_T_2032_en;
  wire [11:0] idxs_T_2035_data;
  wire [5:0] idxs_T_2035_addr;
  wire  idxs_T_2035_en;
  wire [11:0] idxs_T_2038_data;
  wire [5:0] idxs_T_2038_addr;
  wire  idxs_T_2038_en;
  wire [11:0] idxs_T_2041_data;
  wire [5:0] idxs_T_2041_addr;
  wire  idxs_T_2041_en;
  wire [11:0] idxs_T_2044_data;
  wire [5:0] idxs_T_2044_addr;
  wire  idxs_T_2044_en;
  wire [11:0] idxs_T_2047_data;
  wire [5:0] idxs_T_2047_addr;
  wire  idxs_T_2047_en;
  wire [11:0] idxs_T_2050_data;
  wire [5:0] idxs_T_2050_addr;
  wire  idxs_T_2050_en;
  wire [11:0] idxs_T_2053_data;
  wire [5:0] idxs_T_2053_addr;
  wire  idxs_T_2053_en;
  wire [11:0] idxs_T_2056_data;
  wire [5:0] idxs_T_2056_addr;
  wire  idxs_T_2056_en;
  wire [11:0] idxs_T_2059_data;
  wire [5:0] idxs_T_2059_addr;
  wire  idxs_T_2059_en;
  wire [11:0] idxs_T_2062_data;
  wire [5:0] idxs_T_2062_addr;
  wire  idxs_T_2062_en;
  wire [11:0] idxs_T_2065_data;
  wire [5:0] idxs_T_2065_addr;
  wire  idxs_T_2065_en;
  wire [11:0] idxs_T_2068_data;
  wire [5:0] idxs_T_2068_addr;
  wire  idxs_T_2068_en;
  wire [11:0] idxs_T_2071_data;
  wire [5:0] idxs_T_2071_addr;
  wire  idxs_T_2071_en;
  wire [11:0] idxs_T_2074_data;
  wire [5:0] idxs_T_2074_addr;
  wire  idxs_T_2074_en;
  wire [11:0] idxs_T_2077_data;
  wire [5:0] idxs_T_2077_addr;
  wire  idxs_T_2077_en;
  wire [11:0] idxs_T_2080_data;
  wire [5:0] idxs_T_2080_addr;
  wire  idxs_T_2080_en;
  wire [11:0] idxs_T_2083_data;
  wire [5:0] idxs_T_2083_addr;
  wire  idxs_T_2083_en;
  wire [11:0] idxs_T_2086_data;
  wire [5:0] idxs_T_2086_addr;
  wire  idxs_T_2086_en;
  wire [11:0] idxs_T_2089_data;
  wire [5:0] idxs_T_2089_addr;
  wire  idxs_T_2089_en;
  wire [11:0] idxs_T_2092_data;
  wire [5:0] idxs_T_2092_addr;
  wire  idxs_T_2092_en;
  wire [11:0] idxs_T_2095_data;
  wire [5:0] idxs_T_2095_addr;
  wire  idxs_T_2095_en;
  wire [11:0] idxs_T_2098_data;
  wire [5:0] idxs_T_2098_addr;
  wire  idxs_T_2098_en;
  wire [11:0] idxs_T_2101_data;
  wire [5:0] idxs_T_2101_addr;
  wire  idxs_T_2101_en;
  wire [11:0] idxs_T_2104_data;
  wire [5:0] idxs_T_2104_addr;
  wire  idxs_T_2104_en;
  wire [11:0] idxs_T_2107_data;
  wire [5:0] idxs_T_2107_addr;
  wire  idxs_T_2107_en;
  wire [11:0] idxs_T_2110_data;
  wire [5:0] idxs_T_2110_addr;
  wire  idxs_T_2110_en;
  wire [11:0] idxs_T_2113_data;
  wire [5:0] idxs_T_2113_addr;
  wire  idxs_T_2113_en;
  wire [11:0] idxs_T_2116_data;
  wire [5:0] idxs_T_2116_addr;
  wire  idxs_T_2116_en;
  wire [11:0] idxs_T_2119_data;
  wire [5:0] idxs_T_2119_addr;
  wire  idxs_T_2119_en;
  wire [11:0] idxs_T_2122_data;
  wire [5:0] idxs_T_2122_addr;
  wire  idxs_T_2122_en;
  wire [11:0] idxs_T_2125_data;
  wire [5:0] idxs_T_2125_addr;
  wire  idxs_T_2125_en;
  wire [11:0] idxs_T_2128_data;
  wire [5:0] idxs_T_2128_addr;
  wire  idxs_T_2128_en;
  wire [11:0] idxs_T_2131_data;
  wire [5:0] idxs_T_2131_addr;
  wire  idxs_T_2131_en;
  wire [11:0] idxs_T_2134_data;
  wire [5:0] idxs_T_2134_addr;
  wire  idxs_T_2134_en;
  wire [11:0] idxs_T_2137_data;
  wire [5:0] idxs_T_2137_addr;
  wire  idxs_T_2137_en;
  wire [11:0] idxs_T_2140_data;
  wire [5:0] idxs_T_2140_addr;
  wire  idxs_T_2140_en;
  wire [11:0] idxs_T_2143_data;
  wire [5:0] idxs_T_2143_addr;
  wire  idxs_T_2143_en;
  wire [11:0] idxs_T_2146_data;
  wire [5:0] idxs_T_2146_addr;
  wire  idxs_T_2146_en;
  wire [11:0] idxs_T_2149_data;
  wire [5:0] idxs_T_2149_addr;
  wire  idxs_T_2149_en;
  wire [11:0] idxs_T_2152_data;
  wire [5:0] idxs_T_2152_addr;
  wire  idxs_T_2152_en;
  wire [11:0] idxs_T_2155_data;
  wire [5:0] idxs_T_2155_addr;
  wire  idxs_T_2155_en;
  wire [11:0] idxs_T_2872_data;
  wire [5:0] idxs_T_2872_addr;
  wire  idxs_T_2872_mask;
  wire  idxs_T_2872_en;
  reg [2:0] idxPages [0:61];
  reg [31:0] GEN_148;
  wire [2:0] idxPages_T_578_data;
  wire [5:0] idxPages_T_578_addr;
  wire  idxPages_T_578_en;
  wire [2:0] idxPages_T_583_data;
  wire [5:0] idxPages_T_583_addr;
  wire  idxPages_T_583_en;
  wire [2:0] idxPages_T_588_data;
  wire [5:0] idxPages_T_588_addr;
  wire  idxPages_T_588_en;
  wire [2:0] idxPages_T_593_data;
  wire [5:0] idxPages_T_593_addr;
  wire  idxPages_T_593_en;
  wire [2:0] idxPages_T_598_data;
  wire [5:0] idxPages_T_598_addr;
  wire  idxPages_T_598_en;
  wire [2:0] idxPages_T_603_data;
  wire [5:0] idxPages_T_603_addr;
  wire  idxPages_T_603_en;
  wire [2:0] idxPages_T_608_data;
  wire [5:0] idxPages_T_608_addr;
  wire  idxPages_T_608_en;
  wire [2:0] idxPages_T_613_data;
  wire [5:0] idxPages_T_613_addr;
  wire  idxPages_T_613_en;
  wire [2:0] idxPages_T_618_data;
  wire [5:0] idxPages_T_618_addr;
  wire  idxPages_T_618_en;
  wire [2:0] idxPages_T_623_data;
  wire [5:0] idxPages_T_623_addr;
  wire  idxPages_T_623_en;
  wire [2:0] idxPages_T_628_data;
  wire [5:0] idxPages_T_628_addr;
  wire  idxPages_T_628_en;
  wire [2:0] idxPages_T_633_data;
  wire [5:0] idxPages_T_633_addr;
  wire  idxPages_T_633_en;
  wire [2:0] idxPages_T_638_data;
  wire [5:0] idxPages_T_638_addr;
  wire  idxPages_T_638_en;
  wire [2:0] idxPages_T_643_data;
  wire [5:0] idxPages_T_643_addr;
  wire  idxPages_T_643_en;
  wire [2:0] idxPages_T_648_data;
  wire [5:0] idxPages_T_648_addr;
  wire  idxPages_T_648_en;
  wire [2:0] idxPages_T_653_data;
  wire [5:0] idxPages_T_653_addr;
  wire  idxPages_T_653_en;
  wire [2:0] idxPages_T_658_data;
  wire [5:0] idxPages_T_658_addr;
  wire  idxPages_T_658_en;
  wire [2:0] idxPages_T_663_data;
  wire [5:0] idxPages_T_663_addr;
  wire  idxPages_T_663_en;
  wire [2:0] idxPages_T_668_data;
  wire [5:0] idxPages_T_668_addr;
  wire  idxPages_T_668_en;
  wire [2:0] idxPages_T_673_data;
  wire [5:0] idxPages_T_673_addr;
  wire  idxPages_T_673_en;
  wire [2:0] idxPages_T_678_data;
  wire [5:0] idxPages_T_678_addr;
  wire  idxPages_T_678_en;
  wire [2:0] idxPages_T_683_data;
  wire [5:0] idxPages_T_683_addr;
  wire  idxPages_T_683_en;
  wire [2:0] idxPages_T_688_data;
  wire [5:0] idxPages_T_688_addr;
  wire  idxPages_T_688_en;
  wire [2:0] idxPages_T_693_data;
  wire [5:0] idxPages_T_693_addr;
  wire  idxPages_T_693_en;
  wire [2:0] idxPages_T_698_data;
  wire [5:0] idxPages_T_698_addr;
  wire  idxPages_T_698_en;
  wire [2:0] idxPages_T_703_data;
  wire [5:0] idxPages_T_703_addr;
  wire  idxPages_T_703_en;
  wire [2:0] idxPages_T_708_data;
  wire [5:0] idxPages_T_708_addr;
  wire  idxPages_T_708_en;
  wire [2:0] idxPages_T_713_data;
  wire [5:0] idxPages_T_713_addr;
  wire  idxPages_T_713_en;
  wire [2:0] idxPages_T_718_data;
  wire [5:0] idxPages_T_718_addr;
  wire  idxPages_T_718_en;
  wire [2:0] idxPages_T_723_data;
  wire [5:0] idxPages_T_723_addr;
  wire  idxPages_T_723_en;
  wire [2:0] idxPages_T_728_data;
  wire [5:0] idxPages_T_728_addr;
  wire  idxPages_T_728_en;
  wire [2:0] idxPages_T_733_data;
  wire [5:0] idxPages_T_733_addr;
  wire  idxPages_T_733_en;
  wire [2:0] idxPages_T_738_data;
  wire [5:0] idxPages_T_738_addr;
  wire  idxPages_T_738_en;
  wire [2:0] idxPages_T_743_data;
  wire [5:0] idxPages_T_743_addr;
  wire  idxPages_T_743_en;
  wire [2:0] idxPages_T_748_data;
  wire [5:0] idxPages_T_748_addr;
  wire  idxPages_T_748_en;
  wire [2:0] idxPages_T_753_data;
  wire [5:0] idxPages_T_753_addr;
  wire  idxPages_T_753_en;
  wire [2:0] idxPages_T_758_data;
  wire [5:0] idxPages_T_758_addr;
  wire  idxPages_T_758_en;
  wire [2:0] idxPages_T_763_data;
  wire [5:0] idxPages_T_763_addr;
  wire  idxPages_T_763_en;
  wire [2:0] idxPages_T_768_data;
  wire [5:0] idxPages_T_768_addr;
  wire  idxPages_T_768_en;
  wire [2:0] idxPages_T_773_data;
  wire [5:0] idxPages_T_773_addr;
  wire  idxPages_T_773_en;
  wire [2:0] idxPages_T_778_data;
  wire [5:0] idxPages_T_778_addr;
  wire  idxPages_T_778_en;
  wire [2:0] idxPages_T_783_data;
  wire [5:0] idxPages_T_783_addr;
  wire  idxPages_T_783_en;
  wire [2:0] idxPages_T_788_data;
  wire [5:0] idxPages_T_788_addr;
  wire  idxPages_T_788_en;
  wire [2:0] idxPages_T_793_data;
  wire [5:0] idxPages_T_793_addr;
  wire  idxPages_T_793_en;
  wire [2:0] idxPages_T_798_data;
  wire [5:0] idxPages_T_798_addr;
  wire  idxPages_T_798_en;
  wire [2:0] idxPages_T_803_data;
  wire [5:0] idxPages_T_803_addr;
  wire  idxPages_T_803_en;
  wire [2:0] idxPages_T_808_data;
  wire [5:0] idxPages_T_808_addr;
  wire  idxPages_T_808_en;
  wire [2:0] idxPages_T_813_data;
  wire [5:0] idxPages_T_813_addr;
  wire  idxPages_T_813_en;
  wire [2:0] idxPages_T_818_data;
  wire [5:0] idxPages_T_818_addr;
  wire  idxPages_T_818_en;
  wire [2:0] idxPages_T_823_data;
  wire [5:0] idxPages_T_823_addr;
  wire  idxPages_T_823_en;
  wire [2:0] idxPages_T_828_data;
  wire [5:0] idxPages_T_828_addr;
  wire  idxPages_T_828_en;
  wire [2:0] idxPages_T_833_data;
  wire [5:0] idxPages_T_833_addr;
  wire  idxPages_T_833_en;
  wire [2:0] idxPages_T_838_data;
  wire [5:0] idxPages_T_838_addr;
  wire  idxPages_T_838_en;
  wire [2:0] idxPages_T_843_data;
  wire [5:0] idxPages_T_843_addr;
  wire  idxPages_T_843_en;
  wire [2:0] idxPages_T_848_data;
  wire [5:0] idxPages_T_848_addr;
  wire  idxPages_T_848_en;
  wire [2:0] idxPages_T_853_data;
  wire [5:0] idxPages_T_853_addr;
  wire  idxPages_T_853_en;
  wire [2:0] idxPages_T_858_data;
  wire [5:0] idxPages_T_858_addr;
  wire  idxPages_T_858_en;
  wire [2:0] idxPages_T_863_data;
  wire [5:0] idxPages_T_863_addr;
  wire  idxPages_T_863_en;
  wire [2:0] idxPages_T_868_data;
  wire [5:0] idxPages_T_868_addr;
  wire  idxPages_T_868_en;
  wire [2:0] idxPages_T_873_data;
  wire [5:0] idxPages_T_873_addr;
  wire  idxPages_T_873_en;
  wire [2:0] idxPages_T_878_data;
  wire [5:0] idxPages_T_878_addr;
  wire  idxPages_T_878_en;
  wire [2:0] idxPages_T_883_data;
  wire [5:0] idxPages_T_883_addr;
  wire  idxPages_T_883_en;
  wire [2:0] idxPages_T_2874_data;
  wire [5:0] idxPages_T_2874_addr;
  wire  idxPages_T_2874_mask;
  wire  idxPages_T_2874_en;
  reg [11:0] tgts [0:61];
  reg [31:0] GEN_149;
  wire [11:0] tgts_T_3270_data;
  wire [5:0] tgts_T_3270_addr;
  wire  tgts_T_3270_en;
  wire [11:0] tgts_T_3272_data;
  wire [5:0] tgts_T_3272_addr;
  wire  tgts_T_3272_en;
  wire [11:0] tgts_T_3274_data;
  wire [5:0] tgts_T_3274_addr;
  wire  tgts_T_3274_en;
  wire [11:0] tgts_T_3276_data;
  wire [5:0] tgts_T_3276_addr;
  wire  tgts_T_3276_en;
  wire [11:0] tgts_T_3278_data;
  wire [5:0] tgts_T_3278_addr;
  wire  tgts_T_3278_en;
  wire [11:0] tgts_T_3280_data;
  wire [5:0] tgts_T_3280_addr;
  wire  tgts_T_3280_en;
  wire [11:0] tgts_T_3282_data;
  wire [5:0] tgts_T_3282_addr;
  wire  tgts_T_3282_en;
  wire [11:0] tgts_T_3284_data;
  wire [5:0] tgts_T_3284_addr;
  wire  tgts_T_3284_en;
  wire [11:0] tgts_T_3286_data;
  wire [5:0] tgts_T_3286_addr;
  wire  tgts_T_3286_en;
  wire [11:0] tgts_T_3288_data;
  wire [5:0] tgts_T_3288_addr;
  wire  tgts_T_3288_en;
  wire [11:0] tgts_T_3290_data;
  wire [5:0] tgts_T_3290_addr;
  wire  tgts_T_3290_en;
  wire [11:0] tgts_T_3292_data;
  wire [5:0] tgts_T_3292_addr;
  wire  tgts_T_3292_en;
  wire [11:0] tgts_T_3294_data;
  wire [5:0] tgts_T_3294_addr;
  wire  tgts_T_3294_en;
  wire [11:0] tgts_T_3296_data;
  wire [5:0] tgts_T_3296_addr;
  wire  tgts_T_3296_en;
  wire [11:0] tgts_T_3298_data;
  wire [5:0] tgts_T_3298_addr;
  wire  tgts_T_3298_en;
  wire [11:0] tgts_T_3300_data;
  wire [5:0] tgts_T_3300_addr;
  wire  tgts_T_3300_en;
  wire [11:0] tgts_T_3302_data;
  wire [5:0] tgts_T_3302_addr;
  wire  tgts_T_3302_en;
  wire [11:0] tgts_T_3304_data;
  wire [5:0] tgts_T_3304_addr;
  wire  tgts_T_3304_en;
  wire [11:0] tgts_T_3306_data;
  wire [5:0] tgts_T_3306_addr;
  wire  tgts_T_3306_en;
  wire [11:0] tgts_T_3308_data;
  wire [5:0] tgts_T_3308_addr;
  wire  tgts_T_3308_en;
  wire [11:0] tgts_T_3310_data;
  wire [5:0] tgts_T_3310_addr;
  wire  tgts_T_3310_en;
  wire [11:0] tgts_T_3312_data;
  wire [5:0] tgts_T_3312_addr;
  wire  tgts_T_3312_en;
  wire [11:0] tgts_T_3314_data;
  wire [5:0] tgts_T_3314_addr;
  wire  tgts_T_3314_en;
  wire [11:0] tgts_T_3316_data;
  wire [5:0] tgts_T_3316_addr;
  wire  tgts_T_3316_en;
  wire [11:0] tgts_T_3318_data;
  wire [5:0] tgts_T_3318_addr;
  wire  tgts_T_3318_en;
  wire [11:0] tgts_T_3320_data;
  wire [5:0] tgts_T_3320_addr;
  wire  tgts_T_3320_en;
  wire [11:0] tgts_T_3322_data;
  wire [5:0] tgts_T_3322_addr;
  wire  tgts_T_3322_en;
  wire [11:0] tgts_T_3324_data;
  wire [5:0] tgts_T_3324_addr;
  wire  tgts_T_3324_en;
  wire [11:0] tgts_T_3326_data;
  wire [5:0] tgts_T_3326_addr;
  wire  tgts_T_3326_en;
  wire [11:0] tgts_T_3328_data;
  wire [5:0] tgts_T_3328_addr;
  wire  tgts_T_3328_en;
  wire [11:0] tgts_T_3330_data;
  wire [5:0] tgts_T_3330_addr;
  wire  tgts_T_3330_en;
  wire [11:0] tgts_T_3332_data;
  wire [5:0] tgts_T_3332_addr;
  wire  tgts_T_3332_en;
  wire [11:0] tgts_T_3334_data;
  wire [5:0] tgts_T_3334_addr;
  wire  tgts_T_3334_en;
  wire [11:0] tgts_T_3336_data;
  wire [5:0] tgts_T_3336_addr;
  wire  tgts_T_3336_en;
  wire [11:0] tgts_T_3338_data;
  wire [5:0] tgts_T_3338_addr;
  wire  tgts_T_3338_en;
  wire [11:0] tgts_T_3340_data;
  wire [5:0] tgts_T_3340_addr;
  wire  tgts_T_3340_en;
  wire [11:0] tgts_T_3342_data;
  wire [5:0] tgts_T_3342_addr;
  wire  tgts_T_3342_en;
  wire [11:0] tgts_T_3344_data;
  wire [5:0] tgts_T_3344_addr;
  wire  tgts_T_3344_en;
  wire [11:0] tgts_T_3346_data;
  wire [5:0] tgts_T_3346_addr;
  wire  tgts_T_3346_en;
  wire [11:0] tgts_T_3348_data;
  wire [5:0] tgts_T_3348_addr;
  wire  tgts_T_3348_en;
  wire [11:0] tgts_T_3350_data;
  wire [5:0] tgts_T_3350_addr;
  wire  tgts_T_3350_en;
  wire [11:0] tgts_T_3352_data;
  wire [5:0] tgts_T_3352_addr;
  wire  tgts_T_3352_en;
  wire [11:0] tgts_T_3354_data;
  wire [5:0] tgts_T_3354_addr;
  wire  tgts_T_3354_en;
  wire [11:0] tgts_T_3356_data;
  wire [5:0] tgts_T_3356_addr;
  wire  tgts_T_3356_en;
  wire [11:0] tgts_T_3358_data;
  wire [5:0] tgts_T_3358_addr;
  wire  tgts_T_3358_en;
  wire [11:0] tgts_T_3360_data;
  wire [5:0] tgts_T_3360_addr;
  wire  tgts_T_3360_en;
  wire [11:0] tgts_T_3362_data;
  wire [5:0] tgts_T_3362_addr;
  wire  tgts_T_3362_en;
  wire [11:0] tgts_T_3364_data;
  wire [5:0] tgts_T_3364_addr;
  wire  tgts_T_3364_en;
  wire [11:0] tgts_T_3366_data;
  wire [5:0] tgts_T_3366_addr;
  wire  tgts_T_3366_en;
  wire [11:0] tgts_T_3368_data;
  wire [5:0] tgts_T_3368_addr;
  wire  tgts_T_3368_en;
  wire [11:0] tgts_T_3370_data;
  wire [5:0] tgts_T_3370_addr;
  wire  tgts_T_3370_en;
  wire [11:0] tgts_T_3372_data;
  wire [5:0] tgts_T_3372_addr;
  wire  tgts_T_3372_en;
  wire [11:0] tgts_T_3374_data;
  wire [5:0] tgts_T_3374_addr;
  wire  tgts_T_3374_en;
  wire [11:0] tgts_T_3376_data;
  wire [5:0] tgts_T_3376_addr;
  wire  tgts_T_3376_en;
  wire [11:0] tgts_T_3378_data;
  wire [5:0] tgts_T_3378_addr;
  wire  tgts_T_3378_en;
  wire [11:0] tgts_T_3380_data;
  wire [5:0] tgts_T_3380_addr;
  wire  tgts_T_3380_en;
  wire [11:0] tgts_T_3382_data;
  wire [5:0] tgts_T_3382_addr;
  wire  tgts_T_3382_en;
  wire [11:0] tgts_T_3384_data;
  wire [5:0] tgts_T_3384_addr;
  wire  tgts_T_3384_en;
  wire [11:0] tgts_T_3386_data;
  wire [5:0] tgts_T_3386_addr;
  wire  tgts_T_3386_en;
  wire [11:0] tgts_T_3388_data;
  wire [5:0] tgts_T_3388_addr;
  wire  tgts_T_3388_en;
  wire [11:0] tgts_T_3390_data;
  wire [5:0] tgts_T_3390_addr;
  wire  tgts_T_3390_en;
  wire [11:0] tgts_T_3392_data;
  wire [5:0] tgts_T_3392_addr;
  wire  tgts_T_3392_en;
  wire [11:0] tgts_T_2873_data;
  wire [5:0] tgts_T_2873_addr;
  wire  tgts_T_2873_mask;
  wire  tgts_T_2873_en;
  reg [2:0] tgtPages [0:61];
  reg [31:0] GEN_150;
  wire [2:0] tgtPages_T_888_data;
  wire [5:0] tgtPages_T_888_addr;
  wire  tgtPages_T_888_en;
  wire [2:0] tgtPages_T_893_data;
  wire [5:0] tgtPages_T_893_addr;
  wire  tgtPages_T_893_en;
  wire [2:0] tgtPages_T_898_data;
  wire [5:0] tgtPages_T_898_addr;
  wire  tgtPages_T_898_en;
  wire [2:0] tgtPages_T_903_data;
  wire [5:0] tgtPages_T_903_addr;
  wire  tgtPages_T_903_en;
  wire [2:0] tgtPages_T_908_data;
  wire [5:0] tgtPages_T_908_addr;
  wire  tgtPages_T_908_en;
  wire [2:0] tgtPages_T_913_data;
  wire [5:0] tgtPages_T_913_addr;
  wire  tgtPages_T_913_en;
  wire [2:0] tgtPages_T_918_data;
  wire [5:0] tgtPages_T_918_addr;
  wire  tgtPages_T_918_en;
  wire [2:0] tgtPages_T_923_data;
  wire [5:0] tgtPages_T_923_addr;
  wire  tgtPages_T_923_en;
  wire [2:0] tgtPages_T_928_data;
  wire [5:0] tgtPages_T_928_addr;
  wire  tgtPages_T_928_en;
  wire [2:0] tgtPages_T_933_data;
  wire [5:0] tgtPages_T_933_addr;
  wire  tgtPages_T_933_en;
  wire [2:0] tgtPages_T_938_data;
  wire [5:0] tgtPages_T_938_addr;
  wire  tgtPages_T_938_en;
  wire [2:0] tgtPages_T_943_data;
  wire [5:0] tgtPages_T_943_addr;
  wire  tgtPages_T_943_en;
  wire [2:0] tgtPages_T_948_data;
  wire [5:0] tgtPages_T_948_addr;
  wire  tgtPages_T_948_en;
  wire [2:0] tgtPages_T_953_data;
  wire [5:0] tgtPages_T_953_addr;
  wire  tgtPages_T_953_en;
  wire [2:0] tgtPages_T_958_data;
  wire [5:0] tgtPages_T_958_addr;
  wire  tgtPages_T_958_en;
  wire [2:0] tgtPages_T_963_data;
  wire [5:0] tgtPages_T_963_addr;
  wire  tgtPages_T_963_en;
  wire [2:0] tgtPages_T_968_data;
  wire [5:0] tgtPages_T_968_addr;
  wire  tgtPages_T_968_en;
  wire [2:0] tgtPages_T_973_data;
  wire [5:0] tgtPages_T_973_addr;
  wire  tgtPages_T_973_en;
  wire [2:0] tgtPages_T_978_data;
  wire [5:0] tgtPages_T_978_addr;
  wire  tgtPages_T_978_en;
  wire [2:0] tgtPages_T_983_data;
  wire [5:0] tgtPages_T_983_addr;
  wire  tgtPages_T_983_en;
  wire [2:0] tgtPages_T_988_data;
  wire [5:0] tgtPages_T_988_addr;
  wire  tgtPages_T_988_en;
  wire [2:0] tgtPages_T_993_data;
  wire [5:0] tgtPages_T_993_addr;
  wire  tgtPages_T_993_en;
  wire [2:0] tgtPages_T_998_data;
  wire [5:0] tgtPages_T_998_addr;
  wire  tgtPages_T_998_en;
  wire [2:0] tgtPages_T_1003_data;
  wire [5:0] tgtPages_T_1003_addr;
  wire  tgtPages_T_1003_en;
  wire [2:0] tgtPages_T_1008_data;
  wire [5:0] tgtPages_T_1008_addr;
  wire  tgtPages_T_1008_en;
  wire [2:0] tgtPages_T_1013_data;
  wire [5:0] tgtPages_T_1013_addr;
  wire  tgtPages_T_1013_en;
  wire [2:0] tgtPages_T_1018_data;
  wire [5:0] tgtPages_T_1018_addr;
  wire  tgtPages_T_1018_en;
  wire [2:0] tgtPages_T_1023_data;
  wire [5:0] tgtPages_T_1023_addr;
  wire  tgtPages_T_1023_en;
  wire [2:0] tgtPages_T_1028_data;
  wire [5:0] tgtPages_T_1028_addr;
  wire  tgtPages_T_1028_en;
  wire [2:0] tgtPages_T_1033_data;
  wire [5:0] tgtPages_T_1033_addr;
  wire  tgtPages_T_1033_en;
  wire [2:0] tgtPages_T_1038_data;
  wire [5:0] tgtPages_T_1038_addr;
  wire  tgtPages_T_1038_en;
  wire [2:0] tgtPages_T_1043_data;
  wire [5:0] tgtPages_T_1043_addr;
  wire  tgtPages_T_1043_en;
  wire [2:0] tgtPages_T_1048_data;
  wire [5:0] tgtPages_T_1048_addr;
  wire  tgtPages_T_1048_en;
  wire [2:0] tgtPages_T_1053_data;
  wire [5:0] tgtPages_T_1053_addr;
  wire  tgtPages_T_1053_en;
  wire [2:0] tgtPages_T_1058_data;
  wire [5:0] tgtPages_T_1058_addr;
  wire  tgtPages_T_1058_en;
  wire [2:0] tgtPages_T_1063_data;
  wire [5:0] tgtPages_T_1063_addr;
  wire  tgtPages_T_1063_en;
  wire [2:0] tgtPages_T_1068_data;
  wire [5:0] tgtPages_T_1068_addr;
  wire  tgtPages_T_1068_en;
  wire [2:0] tgtPages_T_1073_data;
  wire [5:0] tgtPages_T_1073_addr;
  wire  tgtPages_T_1073_en;
  wire [2:0] tgtPages_T_1078_data;
  wire [5:0] tgtPages_T_1078_addr;
  wire  tgtPages_T_1078_en;
  wire [2:0] tgtPages_T_1083_data;
  wire [5:0] tgtPages_T_1083_addr;
  wire  tgtPages_T_1083_en;
  wire [2:0] tgtPages_T_1088_data;
  wire [5:0] tgtPages_T_1088_addr;
  wire  tgtPages_T_1088_en;
  wire [2:0] tgtPages_T_1093_data;
  wire [5:0] tgtPages_T_1093_addr;
  wire  tgtPages_T_1093_en;
  wire [2:0] tgtPages_T_1098_data;
  wire [5:0] tgtPages_T_1098_addr;
  wire  tgtPages_T_1098_en;
  wire [2:0] tgtPages_T_1103_data;
  wire [5:0] tgtPages_T_1103_addr;
  wire  tgtPages_T_1103_en;
  wire [2:0] tgtPages_T_1108_data;
  wire [5:0] tgtPages_T_1108_addr;
  wire  tgtPages_T_1108_en;
  wire [2:0] tgtPages_T_1113_data;
  wire [5:0] tgtPages_T_1113_addr;
  wire  tgtPages_T_1113_en;
  wire [2:0] tgtPages_T_1118_data;
  wire [5:0] tgtPages_T_1118_addr;
  wire  tgtPages_T_1118_en;
  wire [2:0] tgtPages_T_1123_data;
  wire [5:0] tgtPages_T_1123_addr;
  wire  tgtPages_T_1123_en;
  wire [2:0] tgtPages_T_1128_data;
  wire [5:0] tgtPages_T_1128_addr;
  wire  tgtPages_T_1128_en;
  wire [2:0] tgtPages_T_1133_data;
  wire [5:0] tgtPages_T_1133_addr;
  wire  tgtPages_T_1133_en;
  wire [2:0] tgtPages_T_1138_data;
  wire [5:0] tgtPages_T_1138_addr;
  wire  tgtPages_T_1138_en;
  wire [2:0] tgtPages_T_1143_data;
  wire [5:0] tgtPages_T_1143_addr;
  wire  tgtPages_T_1143_en;
  wire [2:0] tgtPages_T_1148_data;
  wire [5:0] tgtPages_T_1148_addr;
  wire  tgtPages_T_1148_en;
  wire [2:0] tgtPages_T_1153_data;
  wire [5:0] tgtPages_T_1153_addr;
  wire  tgtPages_T_1153_en;
  wire [2:0] tgtPages_T_1158_data;
  wire [5:0] tgtPages_T_1158_addr;
  wire  tgtPages_T_1158_en;
  wire [2:0] tgtPages_T_1163_data;
  wire [5:0] tgtPages_T_1163_addr;
  wire  tgtPages_T_1163_en;
  wire [2:0] tgtPages_T_1168_data;
  wire [5:0] tgtPages_T_1168_addr;
  wire  tgtPages_T_1168_en;
  wire [2:0] tgtPages_T_1173_data;
  wire [5:0] tgtPages_T_1173_addr;
  wire  tgtPages_T_1173_en;
  wire [2:0] tgtPages_T_1178_data;
  wire [5:0] tgtPages_T_1178_addr;
  wire  tgtPages_T_1178_en;
  wire [2:0] tgtPages_T_1183_data;
  wire [5:0] tgtPages_T_1183_addr;
  wire  tgtPages_T_1183_en;
  wire [2:0] tgtPages_T_1188_data;
  wire [5:0] tgtPages_T_1188_addr;
  wire  tgtPages_T_1188_en;
  wire [2:0] tgtPages_T_1193_data;
  wire [5:0] tgtPages_T_1193_addr;
  wire  tgtPages_T_1193_en;
  wire [2:0] tgtPages_T_2875_data;
  wire [5:0] tgtPages_T_2875_addr;
  wire  tgtPages_T_2875_mask;
  wire  tgtPages_T_2875_en;
  reg [26:0] pages [0:5];
  reg [31:0] GEN_151;
  wire [26:0] pages_T_1400_data;
  wire [2:0] pages_T_1400_addr;
  wire  pages_T_1400_en;
  wire [26:0] pages_T_1403_data;
  wire [2:0] pages_T_1403_addr;
  wire  pages_T_1403_en;
  wire [26:0] pages_T_1406_data;
  wire [2:0] pages_T_1406_addr;
  wire  pages_T_1406_en;
  wire [26:0] pages_T_1409_data;
  wire [2:0] pages_T_1409_addr;
  wire  pages_T_1409_en;
  wire [26:0] pages_T_1412_data;
  wire [2:0] pages_T_1412_addr;
  wire  pages_T_1412_en;
  wire [26:0] pages_T_1415_data;
  wire [2:0] pages_T_1415_addr;
  wire  pages_T_1415_en;
  wire [26:0] pages_T_1941_data;
  wire [2:0] pages_T_1941_addr;
  wire  pages_T_1941_en;
  wire [26:0] pages_T_1944_data;
  wire [2:0] pages_T_1944_addr;
  wire  pages_T_1944_en;
  wire [26:0] pages_T_1947_data;
  wire [2:0] pages_T_1947_addr;
  wire  pages_T_1947_en;
  wire [26:0] pages_T_1950_data;
  wire [2:0] pages_T_1950_addr;
  wire  pages_T_1950_en;
  wire [26:0] pages_T_1953_data;
  wire [2:0] pages_T_1953_addr;
  wire  pages_T_1953_en;
  wire [26:0] pages_T_1956_data;
  wire [2:0] pages_T_1956_addr;
  wire  pages_T_1956_en;
  wire [26:0] pages_T_3177_data;
  wire [2:0] pages_T_3177_addr;
  wire  pages_T_3177_en;
  wire [26:0] pages_T_3179_data;
  wire [2:0] pages_T_3179_addr;
  wire  pages_T_3179_en;
  wire [26:0] pages_T_3181_data;
  wire [2:0] pages_T_3181_addr;
  wire  pages_T_3181_en;
  wire [26:0] pages_T_3183_data;
  wire [2:0] pages_T_3183_addr;
  wire  pages_T_3183_en;
  wire [26:0] pages_T_3185_data;
  wire [2:0] pages_T_3185_addr;
  wire  pages_T_3185_en;
  wire [26:0] pages_T_3187_data;
  wire [2:0] pages_T_3187_addr;
  wire  pages_T_3187_en;
  wire [26:0] pages_T_2891_data;
  wire [2:0] pages_T_2891_addr;
  wire  pages_T_2891_mask;
  wire  pages_T_2891_en;
  wire [26:0] pages_T_2895_data;
  wire [2:0] pages_T_2895_addr;
  wire  pages_T_2895_mask;
  wire  pages_T_2895_en;
  wire [26:0] pages_T_2899_data;
  wire [2:0] pages_T_2899_addr;
  wire  pages_T_2899_mask;
  wire  pages_T_2899_en;
  wire [26:0] pages_T_2907_data;
  wire [2:0] pages_T_2907_addr;
  wire  pages_T_2907_mask;
  wire  pages_T_2907_en;
  wire [26:0] pages_T_2911_data;
  wire [2:0] pages_T_2911_addr;
  wire  pages_T_2911_mask;
  wire  pages_T_2911_en;
  wire [26:0] pages_T_2915_data;
  wire [2:0] pages_T_2915_addr;
  wire  pages_T_2915_mask;
  wire  pages_T_2915_en;
  reg [5:0] pageValid;
  reg [31:0] GEN_152;
  wire [7:0] GEN_457;
  wire [7:0] T_580;
  wire [5:0] T_581;
  wire [7:0] T_585;
  wire [5:0] T_586;
  wire [7:0] T_590;
  wire [5:0] T_591;
  wire [7:0] T_595;
  wire [5:0] T_596;
  wire [7:0] T_600;
  wire [5:0] T_601;
  wire [7:0] T_605;
  wire [5:0] T_606;
  wire [7:0] T_610;
  wire [5:0] T_611;
  wire [7:0] T_615;
  wire [5:0] T_616;
  wire [7:0] T_620;
  wire [5:0] T_621;
  wire [7:0] T_625;
  wire [5:0] T_626;
  wire [7:0] T_630;
  wire [5:0] T_631;
  wire [7:0] T_635;
  wire [5:0] T_636;
  wire [7:0] T_640;
  wire [5:0] T_641;
  wire [7:0] T_645;
  wire [5:0] T_646;
  wire [7:0] T_650;
  wire [5:0] T_651;
  wire [7:0] T_655;
  wire [5:0] T_656;
  wire [7:0] T_660;
  wire [5:0] T_661;
  wire [7:0] T_665;
  wire [5:0] T_666;
  wire [7:0] T_670;
  wire [5:0] T_671;
  wire [7:0] T_675;
  wire [5:0] T_676;
  wire [7:0] T_680;
  wire [5:0] T_681;
  wire [7:0] T_685;
  wire [5:0] T_686;
  wire [7:0] T_690;
  wire [5:0] T_691;
  wire [7:0] T_695;
  wire [5:0] T_696;
  wire [7:0] T_700;
  wire [5:0] T_701;
  wire [7:0] T_705;
  wire [5:0] T_706;
  wire [7:0] T_710;
  wire [5:0] T_711;
  wire [7:0] T_715;
  wire [5:0] T_716;
  wire [7:0] T_720;
  wire [5:0] T_721;
  wire [7:0] T_725;
  wire [5:0] T_726;
  wire [7:0] T_730;
  wire [5:0] T_731;
  wire [7:0] T_735;
  wire [5:0] T_736;
  wire [7:0] T_740;
  wire [5:0] T_741;
  wire [7:0] T_745;
  wire [5:0] T_746;
  wire [7:0] T_750;
  wire [5:0] T_751;
  wire [7:0] T_755;
  wire [5:0] T_756;
  wire [7:0] T_760;
  wire [5:0] T_761;
  wire [7:0] T_765;
  wire [5:0] T_766;
  wire [7:0] T_770;
  wire [5:0] T_771;
  wire [7:0] T_775;
  wire [5:0] T_776;
  wire [7:0] T_780;
  wire [5:0] T_781;
  wire [7:0] T_785;
  wire [5:0] T_786;
  wire [7:0] T_790;
  wire [5:0] T_791;
  wire [7:0] T_795;
  wire [5:0] T_796;
  wire [7:0] T_800;
  wire [5:0] T_801;
  wire [7:0] T_805;
  wire [5:0] T_806;
  wire [7:0] T_810;
  wire [5:0] T_811;
  wire [7:0] T_815;
  wire [5:0] T_816;
  wire [7:0] T_820;
  wire [5:0] T_821;
  wire [7:0] T_825;
  wire [5:0] T_826;
  wire [7:0] T_830;
  wire [5:0] T_831;
  wire [7:0] T_835;
  wire [5:0] T_836;
  wire [7:0] T_840;
  wire [5:0] T_841;
  wire [7:0] T_845;
  wire [5:0] T_846;
  wire [7:0] T_850;
  wire [5:0] T_851;
  wire [7:0] T_855;
  wire [5:0] T_856;
  wire [7:0] T_860;
  wire [5:0] T_861;
  wire [7:0] T_865;
  wire [5:0] T_866;
  wire [7:0] T_870;
  wire [5:0] T_871;
  wire [7:0] T_875;
  wire [5:0] T_876;
  wire [7:0] T_880;
  wire [5:0] T_881;
  wire [7:0] T_885;
  wire [5:0] T_886;
  wire [7:0] T_890;
  wire [5:0] T_891;
  wire [7:0] T_895;
  wire [5:0] T_896;
  wire [7:0] T_900;
  wire [5:0] T_901;
  wire [7:0] T_905;
  wire [5:0] T_906;
  wire [7:0] T_910;
  wire [5:0] T_911;
  wire [7:0] T_915;
  wire [5:0] T_916;
  wire [7:0] T_920;
  wire [5:0] T_921;
  wire [7:0] T_925;
  wire [5:0] T_926;
  wire [7:0] T_930;
  wire [5:0] T_931;
  wire [7:0] T_935;
  wire [5:0] T_936;
  wire [7:0] T_940;
  wire [5:0] T_941;
  wire [7:0] T_945;
  wire [5:0] T_946;
  wire [7:0] T_950;
  wire [5:0] T_951;
  wire [7:0] T_955;
  wire [5:0] T_956;
  wire [7:0] T_960;
  wire [5:0] T_961;
  wire [7:0] T_965;
  wire [5:0] T_966;
  wire [7:0] T_970;
  wire [5:0] T_971;
  wire [7:0] T_975;
  wire [5:0] T_976;
  wire [7:0] T_980;
  wire [5:0] T_981;
  wire [7:0] T_985;
  wire [5:0] T_986;
  wire [7:0] T_990;
  wire [5:0] T_991;
  wire [7:0] T_995;
  wire [5:0] T_996;
  wire [7:0] T_1000;
  wire [5:0] T_1001;
  wire [7:0] T_1005;
  wire [5:0] T_1006;
  wire [7:0] T_1010;
  wire [5:0] T_1011;
  wire [7:0] T_1015;
  wire [5:0] T_1016;
  wire [7:0] T_1020;
  wire [5:0] T_1021;
  wire [7:0] T_1025;
  wire [5:0] T_1026;
  wire [7:0] T_1030;
  wire [5:0] T_1031;
  wire [7:0] T_1035;
  wire [5:0] T_1036;
  wire [7:0] T_1040;
  wire [5:0] T_1041;
  wire [7:0] T_1045;
  wire [5:0] T_1046;
  wire [7:0] T_1050;
  wire [5:0] T_1051;
  wire [7:0] T_1055;
  wire [5:0] T_1056;
  wire [7:0] T_1060;
  wire [5:0] T_1061;
  wire [7:0] T_1065;
  wire [5:0] T_1066;
  wire [7:0] T_1070;
  wire [5:0] T_1071;
  wire [7:0] T_1075;
  wire [5:0] T_1076;
  wire [7:0] T_1080;
  wire [5:0] T_1081;
  wire [7:0] T_1085;
  wire [5:0] T_1086;
  wire [7:0] T_1090;
  wire [5:0] T_1091;
  wire [7:0] T_1095;
  wire [5:0] T_1096;
  wire [7:0] T_1100;
  wire [5:0] T_1101;
  wire [7:0] T_1105;
  wire [5:0] T_1106;
  wire [7:0] T_1110;
  wire [5:0] T_1111;
  wire [7:0] T_1115;
  wire [5:0] T_1116;
  wire [7:0] T_1120;
  wire [5:0] T_1121;
  wire [7:0] T_1125;
  wire [5:0] T_1126;
  wire [7:0] T_1130;
  wire [5:0] T_1131;
  wire [7:0] T_1135;
  wire [5:0] T_1136;
  wire [7:0] T_1140;
  wire [5:0] T_1141;
  wire [7:0] T_1145;
  wire [5:0] T_1146;
  wire [7:0] T_1150;
  wire [5:0] T_1151;
  wire [7:0] T_1155;
  wire [5:0] T_1156;
  wire [7:0] T_1160;
  wire [5:0] T_1161;
  wire [7:0] T_1165;
  wire [5:0] T_1166;
  wire [7:0] T_1170;
  wire [5:0] T_1171;
  wire [7:0] T_1175;
  wire [5:0] T_1176;
  wire [7:0] T_1180;
  wire [5:0] T_1181;
  wire [7:0] T_1185;
  wire [5:0] T_1186;
  wire [7:0] T_1190;
  wire [5:0] T_1191;
  wire [7:0] T_1195;
  wire [5:0] T_1196;
  reg  useRAS_0;
  reg [31:0] GEN_153;
  reg  useRAS_1;
  reg [31:0] GEN_154;
  reg  useRAS_2;
  reg [31:0] GEN_155;
  reg  useRAS_3;
  reg [31:0] GEN_156;
  reg  useRAS_4;
  reg [31:0] GEN_157;
  reg  useRAS_5;
  reg [31:0] GEN_158;
  reg  useRAS_6;
  reg [31:0] GEN_159;
  reg  useRAS_7;
  reg [31:0] GEN_160;
  reg  useRAS_8;
  reg [31:0] GEN_161;
  reg  useRAS_9;
  reg [31:0] GEN_162;
  reg  useRAS_10;
  reg [31:0] GEN_163;
  reg  useRAS_11;
  reg [31:0] GEN_164;
  reg  useRAS_12;
  reg [31:0] GEN_165;
  reg  useRAS_13;
  reg [31:0] GEN_166;
  reg  useRAS_14;
  reg [31:0] GEN_167;
  reg  useRAS_15;
  reg [31:0] GEN_168;
  reg  useRAS_16;
  reg [31:0] GEN_169;
  reg  useRAS_17;
  reg [31:0] GEN_170;
  reg  useRAS_18;
  reg [31:0] GEN_171;
  reg  useRAS_19;
  reg [31:0] GEN_172;
  reg  useRAS_20;
  reg [31:0] GEN_173;
  reg  useRAS_21;
  reg [31:0] GEN_174;
  reg  useRAS_22;
  reg [31:0] GEN_175;
  reg  useRAS_23;
  reg [31:0] GEN_177;
  reg  useRAS_24;
  reg [31:0] GEN_178;
  reg  useRAS_25;
  reg [31:0] GEN_179;
  reg  useRAS_26;
  reg [31:0] GEN_180;
  reg  useRAS_27;
  reg [31:0] GEN_181;
  reg  useRAS_28;
  reg [31:0] GEN_182;
  reg  useRAS_29;
  reg [31:0] GEN_183;
  reg  useRAS_30;
  reg [31:0] GEN_184;
  reg  useRAS_31;
  reg [31:0] GEN_185;
  reg  useRAS_32;
  reg [31:0] GEN_186;
  reg  useRAS_33;
  reg [31:0] GEN_187;
  reg  useRAS_34;
  reg [31:0] GEN_188;
  reg  useRAS_35;
  reg [31:0] GEN_189;
  reg  useRAS_36;
  reg [31:0] GEN_190;
  reg  useRAS_37;
  reg [31:0] GEN_191;
  reg  useRAS_38;
  reg [31:0] GEN_192;
  reg  useRAS_39;
  reg [31:0] GEN_193;
  reg  useRAS_40;
  reg [31:0] GEN_194;
  reg  useRAS_41;
  reg [31:0] GEN_195;
  reg  useRAS_42;
  reg [31:0] GEN_196;
  reg  useRAS_43;
  reg [31:0] GEN_197;
  reg  useRAS_44;
  reg [31:0] GEN_198;
  reg  useRAS_45;
  reg [31:0] GEN_199;
  reg  useRAS_46;
  reg [31:0] GEN_200;
  reg  useRAS_47;
  reg [31:0] GEN_201;
  reg  useRAS_48;
  reg [31:0] GEN_202;
  reg  useRAS_49;
  reg [31:0] GEN_203;
  reg  useRAS_50;
  reg [31:0] GEN_204;
  reg  useRAS_51;
  reg [31:0] GEN_205;
  reg  useRAS_52;
  reg [31:0] GEN_206;
  reg  useRAS_53;
  reg [31:0] GEN_207;
  reg  useRAS_54;
  reg [31:0] GEN_208;
  reg  useRAS_55;
  reg [31:0] GEN_209;
  reg  useRAS_56;
  reg [31:0] GEN_210;
  reg  useRAS_57;
  reg [31:0] GEN_211;
  reg  useRAS_58;
  reg [31:0] GEN_212;
  reg  useRAS_59;
  reg [31:0] GEN_213;
  reg  useRAS_60;
  reg [31:0] GEN_214;
  reg  useRAS_61;
  reg [31:0] GEN_215;
  reg  isJump_0;
  reg [31:0] GEN_216;
  reg  isJump_1;
  reg [31:0] GEN_217;
  reg  isJump_2;
  reg [31:0] GEN_218;
  reg  isJump_3;
  reg [31:0] GEN_219;
  reg  isJump_4;
  reg [31:0] GEN_220;
  reg  isJump_5;
  reg [31:0] GEN_221;
  reg  isJump_6;
  reg [31:0] GEN_222;
  reg  isJump_7;
  reg [31:0] GEN_223;
  reg  isJump_8;
  reg [31:0] GEN_224;
  reg  isJump_9;
  reg [31:0] GEN_225;
  reg  isJump_10;
  reg [31:0] GEN_226;
  reg  isJump_11;
  reg [31:0] GEN_227;
  reg  isJump_12;
  reg [31:0] GEN_228;
  reg  isJump_13;
  reg [31:0] GEN_229;
  reg  isJump_14;
  reg [31:0] GEN_230;
  reg  isJump_15;
  reg [31:0] GEN_231;
  reg  isJump_16;
  reg [31:0] GEN_232;
  reg  isJump_17;
  reg [31:0] GEN_233;
  reg  isJump_18;
  reg [31:0] GEN_234;
  reg  isJump_19;
  reg [31:0] GEN_235;
  reg  isJump_20;
  reg [31:0] GEN_236;
  reg  isJump_21;
  reg [31:0] GEN_237;
  reg  isJump_22;
  reg [31:0] GEN_238;
  reg  isJump_23;
  reg [31:0] GEN_240;
  reg  isJump_24;
  reg [31:0] GEN_241;
  reg  isJump_25;
  reg [31:0] GEN_242;
  reg  isJump_26;
  reg [31:0] GEN_243;
  reg  isJump_27;
  reg [31:0] GEN_244;
  reg  isJump_28;
  reg [31:0] GEN_245;
  reg  isJump_29;
  reg [31:0] GEN_246;
  reg  isJump_30;
  reg [31:0] GEN_247;
  reg  isJump_31;
  reg [31:0] GEN_248;
  reg  isJump_32;
  reg [31:0] GEN_249;
  reg  isJump_33;
  reg [31:0] GEN_250;
  reg  isJump_34;
  reg [31:0] GEN_251;
  reg  isJump_35;
  reg [31:0] GEN_252;
  reg  isJump_36;
  reg [31:0] GEN_253;
  reg  isJump_37;
  reg [31:0] GEN_254;
  reg  isJump_38;
  reg [31:0] GEN_255;
  reg  isJump_39;
  reg [31:0] GEN_256;
  reg  isJump_40;
  reg [31:0] GEN_257;
  reg  isJump_41;
  reg [31:0] GEN_258;
  reg  isJump_42;
  reg [31:0] GEN_259;
  reg  isJump_43;
  reg [31:0] GEN_260;
  reg  isJump_44;
  reg [31:0] GEN_323;
  reg  isJump_45;
  reg [31:0] GEN_386;
  reg  isJump_46;
  reg [31:0] GEN_387;
  reg  isJump_47;
  reg [31:0] GEN_388;
  reg  isJump_48;
  reg [31:0] GEN_389;
  reg  isJump_49;
  reg [31:0] GEN_390;
  reg  isJump_50;
  reg [31:0] GEN_391;
  reg  isJump_51;
  reg [31:0] GEN_392;
  reg  isJump_52;
  reg [31:0] GEN_394;
  reg  isJump_53;
  reg [31:0] GEN_395;
  reg  isJump_54;
  reg [31:0] GEN_396;
  reg  isJump_55;
  reg [31:0] GEN_397;
  reg  isJump_56;
  reg [31:0] GEN_399;
  reg  isJump_57;
  reg [31:0] GEN_400;
  reg  isJump_58;
  reg [31:0] GEN_401;
  reg  isJump_59;
  reg [31:0] GEN_402;
  reg  isJump_60;
  reg [31:0] GEN_404;
  reg  isJump_61;
  reg [31:0] GEN_405;
  reg  brIdx [0:61];
  reg [31:0] GEN_406;
  wire  brIdx_T_3612_data;
  wire [5:0] brIdx_T_3612_addr;
  wire  brIdx_T_3612_en;
  wire  brIdx_T_2876_data;
  wire [5:0] brIdx_T_2876_addr;
  wire  brIdx_T_2876_mask;
  wire  brIdx_T_2876_en;
  reg  T_1215;
  reg [31:0] GEN_407;
  reg  T_1216_prediction_valid;
  reg [31:0] GEN_409;
  reg  T_1216_prediction_bits_taken;
  reg [31:0] GEN_410;
  reg  T_1216_prediction_bits_mask;
  reg [31:0] GEN_411;
  reg  T_1216_prediction_bits_bridx;
  reg [31:0] GEN_412;
  reg [38:0] T_1216_prediction_bits_target;
  reg [63:0] GEN_414;
  reg [5:0] T_1216_prediction_bits_entry;
  reg [31:0] GEN_415;
  reg [6:0] T_1216_prediction_bits_bht_history;
  reg [31:0] GEN_416;
  reg [1:0] T_1216_prediction_bits_bht_value;
  reg [31:0] GEN_417;
  reg [38:0] T_1216_pc;
  reg [63:0] GEN_419;
  reg [38:0] T_1216_target;
  reg [63:0] GEN_420;
  reg  T_1216_taken;
  reg [31:0] GEN_426;
  reg  T_1216_isJump;
  reg [31:0] GEN_427;
  reg  T_1216_isReturn;
  reg [31:0] GEN_428;
  reg [38:0] T_1216_br_pc;
  reg [63:0] GEN_429;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [38:0] GEN_8;
  wire [5:0] GEN_9;
  wire [6:0] GEN_10;
  wire [1:0] GEN_11;
  wire [38:0] GEN_12;
  wire [38:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [38:0] GEN_17;
  wire  r_btb_update_valid;
  wire  r_btb_update_bits_prediction_valid;
  wire  r_btb_update_bits_prediction_bits_taken;
  wire  r_btb_update_bits_prediction_bits_mask;
  wire  r_btb_update_bits_prediction_bits_bridx;
  wire [38:0] r_btb_update_bits_prediction_bits_target;
  wire [5:0] r_btb_update_bits_prediction_bits_entry;
  wire [6:0] r_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] r_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] r_btb_update_bits_pc;
  wire [38:0] r_btb_update_bits_target;
  wire  r_btb_update_bits_taken;
  wire  r_btb_update_bits_isJump;
  wire  r_btb_update_bits_isReturn;
  wire [38:0] r_btb_update_bits_br_pc;
  wire [26:0] T_1398;
  wire  T_1401;
  wire  T_1404;
  wire  T_1407;
  wire  T_1410;
  wire  T_1413;
  wire  T_1416;
  wire  T_1422_0;
  wire  T_1422_1;
  wire  T_1422_2;
  wire  T_1422_3;
  wire  T_1422_4;
  wire  T_1422_5;
  wire [1:0] T_1424;
  wire [2:0] T_1425;
  wire [1:0] T_1426;
  wire [2:0] T_1427;
  wire [5:0] T_1428;
  wire [5:0] pageHit;
  wire [11:0] T_1429;
  wire  T_1432;
  wire  T_1435;
  wire  T_1438;
  wire  T_1441;
  wire  T_1444;
  wire  T_1447;
  wire  T_1450;
  wire  T_1453;
  wire  T_1456;
  wire  T_1459;
  wire  T_1462;
  wire  T_1465;
  wire  T_1468;
  wire  T_1471;
  wire  T_1474;
  wire  T_1477;
  wire  T_1480;
  wire  T_1483;
  wire  T_1486;
  wire  T_1489;
  wire  T_1492;
  wire  T_1495;
  wire  T_1498;
  wire  T_1501;
  wire  T_1504;
  wire  T_1507;
  wire  T_1510;
  wire  T_1513;
  wire  T_1516;
  wire  T_1519;
  wire  T_1522;
  wire  T_1525;
  wire  T_1528;
  wire  T_1531;
  wire  T_1534;
  wire  T_1537;
  wire  T_1540;
  wire  T_1543;
  wire  T_1546;
  wire  T_1549;
  wire  T_1552;
  wire  T_1555;
  wire  T_1558;
  wire  T_1561;
  wire  T_1564;
  wire  T_1567;
  wire  T_1570;
  wire  T_1573;
  wire  T_1576;
  wire  T_1579;
  wire  T_1582;
  wire  T_1585;
  wire  T_1588;
  wire  T_1591;
  wire  T_1594;
  wire  T_1597;
  wire  T_1600;
  wire  T_1603;
  wire  T_1606;
  wire  T_1609;
  wire  T_1612;
  wire  T_1615;
  wire  T_1621_0;
  wire  T_1621_1;
  wire  T_1621_2;
  wire  T_1621_3;
  wire  T_1621_4;
  wire  T_1621_5;
  wire  T_1621_6;
  wire  T_1621_7;
  wire  T_1621_8;
  wire  T_1621_9;
  wire  T_1621_10;
  wire  T_1621_11;
  wire  T_1621_12;
  wire  T_1621_13;
  wire  T_1621_14;
  wire  T_1621_15;
  wire  T_1621_16;
  wire  T_1621_17;
  wire  T_1621_18;
  wire  T_1621_19;
  wire  T_1621_20;
  wire  T_1621_21;
  wire  T_1621_22;
  wire  T_1621_23;
  wire  T_1621_24;
  wire  T_1621_25;
  wire  T_1621_26;
  wire  T_1621_27;
  wire  T_1621_28;
  wire  T_1621_29;
  wire  T_1621_30;
  wire  T_1621_31;
  wire  T_1621_32;
  wire  T_1621_33;
  wire  T_1621_34;
  wire  T_1621_35;
  wire  T_1621_36;
  wire  T_1621_37;
  wire  T_1621_38;
  wire  T_1621_39;
  wire  T_1621_40;
  wire  T_1621_41;
  wire  T_1621_42;
  wire  T_1621_43;
  wire  T_1621_44;
  wire  T_1621_45;
  wire  T_1621_46;
  wire  T_1621_47;
  wire  T_1621_48;
  wire  T_1621_49;
  wire  T_1621_50;
  wire  T_1621_51;
  wire  T_1621_52;
  wire  T_1621_53;
  wire  T_1621_54;
  wire  T_1621_55;
  wire  T_1621_56;
  wire  T_1621_57;
  wire  T_1621_58;
  wire  T_1621_59;
  wire  T_1621_60;
  wire  T_1621_61;
  wire [1:0] T_1623;
  wire [2:0] T_1624;
  wire [1:0] T_1625;
  wire [1:0] T_1626;
  wire [3:0] T_1627;
  wire [6:0] T_1628;
  wire [1:0] T_1629;
  wire [1:0] T_1630;
  wire [3:0] T_1631;
  wire [1:0] T_1632;
  wire [1:0] T_1633;
  wire [3:0] T_1634;
  wire [7:0] T_1635;
  wire [14:0] T_1636;
  wire [1:0] T_1637;
  wire [1:0] T_1638;
  wire [3:0] T_1639;
  wire [1:0] T_1640;
  wire [1:0] T_1641;
  wire [3:0] T_1642;
  wire [7:0] T_1643;
  wire [1:0] T_1644;
  wire [1:0] T_1645;
  wire [3:0] T_1646;
  wire [1:0] T_1647;
  wire [1:0] T_1648;
  wire [3:0] T_1649;
  wire [7:0] T_1650;
  wire [15:0] T_1651;
  wire [30:0] T_1652;
  wire [1:0] T_1653;
  wire [2:0] T_1654;
  wire [1:0] T_1655;
  wire [1:0] T_1656;
  wire [3:0] T_1657;
  wire [6:0] T_1658;
  wire [1:0] T_1659;
  wire [1:0] T_1660;
  wire [3:0] T_1661;
  wire [1:0] T_1662;
  wire [1:0] T_1663;
  wire [3:0] T_1664;
  wire [7:0] T_1665;
  wire [14:0] T_1666;
  wire [1:0] T_1667;
  wire [1:0] T_1668;
  wire [3:0] T_1669;
  wire [1:0] T_1670;
  wire [1:0] T_1671;
  wire [3:0] T_1672;
  wire [7:0] T_1673;
  wire [1:0] T_1674;
  wire [1:0] T_1675;
  wire [3:0] T_1676;
  wire [1:0] T_1677;
  wire [1:0] T_1678;
  wire [3:0] T_1679;
  wire [7:0] T_1680;
  wire [15:0] T_1681;
  wire [30:0] T_1682;
  wire [61:0] T_1683;
  wire [5:0] T_1684;
  wire [5:0] T_1685;
  wire [5:0] T_1686;
  wire [5:0] T_1687;
  wire [5:0] T_1688;
  wire [5:0] T_1689;
  wire [5:0] T_1690;
  wire [5:0] T_1691;
  wire [5:0] T_1692;
  wire [5:0] T_1693;
  wire [5:0] T_1694;
  wire [5:0] T_1695;
  wire [5:0] T_1696;
  wire [5:0] T_1697;
  wire [5:0] T_1698;
  wire [5:0] T_1699;
  wire [5:0] T_1700;
  wire [5:0] T_1701;
  wire [5:0] T_1702;
  wire [5:0] T_1703;
  wire [5:0] T_1704;
  wire [5:0] T_1705;
  wire [5:0] T_1706;
  wire [5:0] T_1707;
  wire [5:0] T_1708;
  wire [5:0] T_1709;
  wire [5:0] T_1710;
  wire [5:0] T_1711;
  wire [5:0] T_1712;
  wire [5:0] T_1713;
  wire [5:0] T_1714;
  wire [5:0] T_1715;
  wire [5:0] T_1716;
  wire [5:0] T_1717;
  wire [5:0] T_1718;
  wire [5:0] T_1719;
  wire [5:0] T_1720;
  wire [5:0] T_1721;
  wire [5:0] T_1722;
  wire [5:0] T_1723;
  wire [5:0] T_1724;
  wire [5:0] T_1725;
  wire [5:0] T_1726;
  wire [5:0] T_1727;
  wire [5:0] T_1728;
  wire [5:0] T_1729;
  wire [5:0] T_1730;
  wire [5:0] T_1731;
  wire [5:0] T_1732;
  wire [5:0] T_1733;
  wire [5:0] T_1734;
  wire [5:0] T_1735;
  wire [5:0] T_1736;
  wire [5:0] T_1737;
  wire [5:0] T_1738;
  wire [5:0] T_1739;
  wire [5:0] T_1740;
  wire [5:0] T_1741;
  wire [5:0] T_1742;
  wire [5:0] T_1743;
  wire [5:0] T_1744;
  wire [5:0] T_1745;
  wire [5:0] GEN_581;
  wire  T_1747;
  wire  T_1749;
  wire  T_1751;
  wire  T_1753;
  wire  T_1755;
  wire  T_1757;
  wire  T_1759;
  wire  T_1761;
  wire  T_1763;
  wire  T_1765;
  wire  T_1767;
  wire  T_1769;
  wire  T_1771;
  wire  T_1773;
  wire  T_1775;
  wire  T_1777;
  wire  T_1779;
  wire  T_1781;
  wire  T_1783;
  wire  T_1785;
  wire  T_1787;
  wire  T_1789;
  wire  T_1791;
  wire  T_1793;
  wire  T_1795;
  wire  T_1797;
  wire  T_1799;
  wire  T_1801;
  wire  T_1803;
  wire  T_1805;
  wire  T_1807;
  wire  T_1809;
  wire  T_1811;
  wire  T_1813;
  wire  T_1815;
  wire  T_1817;
  wire  T_1819;
  wire  T_1821;
  wire  T_1823;
  wire  T_1825;
  wire  T_1827;
  wire  T_1829;
  wire  T_1831;
  wire  T_1833;
  wire  T_1835;
  wire  T_1837;
  wire  T_1839;
  wire  T_1841;
  wire  T_1843;
  wire  T_1845;
  wire  T_1847;
  wire  T_1849;
  wire  T_1851;
  wire  T_1853;
  wire  T_1855;
  wire  T_1857;
  wire  T_1859;
  wire  T_1861;
  wire  T_1863;
  wire  T_1865;
  wire  T_1867;
  wire  T_1869;
  wire  T_1875_0;
  wire  T_1875_1;
  wire  T_1875_2;
  wire  T_1875_3;
  wire  T_1875_4;
  wire  T_1875_5;
  wire  T_1875_6;
  wire  T_1875_7;
  wire  T_1875_8;
  wire  T_1875_9;
  wire  T_1875_10;
  wire  T_1875_11;
  wire  T_1875_12;
  wire  T_1875_13;
  wire  T_1875_14;
  wire  T_1875_15;
  wire  T_1875_16;
  wire  T_1875_17;
  wire  T_1875_18;
  wire  T_1875_19;
  wire  T_1875_20;
  wire  T_1875_21;
  wire  T_1875_22;
  wire  T_1875_23;
  wire  T_1875_24;
  wire  T_1875_25;
  wire  T_1875_26;
  wire  T_1875_27;
  wire  T_1875_28;
  wire  T_1875_29;
  wire  T_1875_30;
  wire  T_1875_31;
  wire  T_1875_32;
  wire  T_1875_33;
  wire  T_1875_34;
  wire  T_1875_35;
  wire  T_1875_36;
  wire  T_1875_37;
  wire  T_1875_38;
  wire  T_1875_39;
  wire  T_1875_40;
  wire  T_1875_41;
  wire  T_1875_42;
  wire  T_1875_43;
  wire  T_1875_44;
  wire  T_1875_45;
  wire  T_1875_46;
  wire  T_1875_47;
  wire  T_1875_48;
  wire  T_1875_49;
  wire  T_1875_50;
  wire  T_1875_51;
  wire  T_1875_52;
  wire  T_1875_53;
  wire  T_1875_54;
  wire  T_1875_55;
  wire  T_1875_56;
  wire  T_1875_57;
  wire  T_1875_58;
  wire  T_1875_59;
  wire  T_1875_60;
  wire  T_1875_61;
  wire [1:0] T_1877;
  wire [2:0] T_1878;
  wire [1:0] T_1879;
  wire [1:0] T_1880;
  wire [3:0] T_1881;
  wire [6:0] T_1882;
  wire [1:0] T_1883;
  wire [1:0] T_1884;
  wire [3:0] T_1885;
  wire [1:0] T_1886;
  wire [1:0] T_1887;
  wire [3:0] T_1888;
  wire [7:0] T_1889;
  wire [14:0] T_1890;
  wire [1:0] T_1891;
  wire [1:0] T_1892;
  wire [3:0] T_1893;
  wire [1:0] T_1894;
  wire [1:0] T_1895;
  wire [3:0] T_1896;
  wire [7:0] T_1897;
  wire [1:0] T_1898;
  wire [1:0] T_1899;
  wire [3:0] T_1900;
  wire [1:0] T_1901;
  wire [1:0] T_1902;
  wire [3:0] T_1903;
  wire [7:0] T_1904;
  wire [15:0] T_1905;
  wire [30:0] T_1906;
  wire [1:0] T_1907;
  wire [2:0] T_1908;
  wire [1:0] T_1909;
  wire [1:0] T_1910;
  wire [3:0] T_1911;
  wire [6:0] T_1912;
  wire [1:0] T_1913;
  wire [1:0] T_1914;
  wire [3:0] T_1915;
  wire [1:0] T_1916;
  wire [1:0] T_1917;
  wire [3:0] T_1918;
  wire [7:0] T_1919;
  wire [14:0] T_1920;
  wire [1:0] T_1921;
  wire [1:0] T_1922;
  wire [3:0] T_1923;
  wire [1:0] T_1924;
  wire [1:0] T_1925;
  wire [3:0] T_1926;
  wire [7:0] T_1927;
  wire [1:0] T_1928;
  wire [1:0] T_1929;
  wire [3:0] T_1930;
  wire [1:0] T_1931;
  wire [1:0] T_1932;
  wire [3:0] T_1933;
  wire [7:0] T_1934;
  wire [15:0] T_1935;
  wire [30:0] T_1936;
  wire [61:0] T_1937;
  wire [61:0] T_1938;
  wire [61:0] hits;
  wire [26:0] T_1939;
  wire  T_1942;
  wire  T_1945;
  wire  T_1948;
  wire  T_1951;
  wire  T_1954;
  wire  T_1957;
  wire  T_1963_0;
  wire  T_1963_1;
  wire  T_1963_2;
  wire  T_1963_3;
  wire  T_1963_4;
  wire  T_1963_5;
  wire [1:0] T_1965;
  wire [2:0] T_1966;
  wire [1:0] T_1967;
  wire [2:0] T_1968;
  wire [5:0] T_1969;
  wire [5:0] updatePageHit;
  wire [11:0] T_1970;
  wire  T_1973;
  wire  T_1976;
  wire  T_1979;
  wire  T_1982;
  wire  T_1985;
  wire  T_1988;
  wire  T_1991;
  wire  T_1994;
  wire  T_1997;
  wire  T_2000;
  wire  T_2003;
  wire  T_2006;
  wire  T_2009;
  wire  T_2012;
  wire  T_2015;
  wire  T_2018;
  wire  T_2021;
  wire  T_2024;
  wire  T_2027;
  wire  T_2030;
  wire  T_2033;
  wire  T_2036;
  wire  T_2039;
  wire  T_2042;
  wire  T_2045;
  wire  T_2048;
  wire  T_2051;
  wire  T_2054;
  wire  T_2057;
  wire  T_2060;
  wire  T_2063;
  wire  T_2066;
  wire  T_2069;
  wire  T_2072;
  wire  T_2075;
  wire  T_2078;
  wire  T_2081;
  wire  T_2084;
  wire  T_2087;
  wire  T_2090;
  wire  T_2093;
  wire  T_2096;
  wire  T_2099;
  wire  T_2102;
  wire  T_2105;
  wire  T_2108;
  wire  T_2111;
  wire  T_2114;
  wire  T_2117;
  wire  T_2120;
  wire  T_2123;
  wire  T_2126;
  wire  T_2129;
  wire  T_2132;
  wire  T_2135;
  wire  T_2138;
  wire  T_2141;
  wire  T_2144;
  wire  T_2147;
  wire  T_2150;
  wire  T_2153;
  wire  T_2156;
  wire  T_2162_0;
  wire  T_2162_1;
  wire  T_2162_2;
  wire  T_2162_3;
  wire  T_2162_4;
  wire  T_2162_5;
  wire  T_2162_6;
  wire  T_2162_7;
  wire  T_2162_8;
  wire  T_2162_9;
  wire  T_2162_10;
  wire  T_2162_11;
  wire  T_2162_12;
  wire  T_2162_13;
  wire  T_2162_14;
  wire  T_2162_15;
  wire  T_2162_16;
  wire  T_2162_17;
  wire  T_2162_18;
  wire  T_2162_19;
  wire  T_2162_20;
  wire  T_2162_21;
  wire  T_2162_22;
  wire  T_2162_23;
  wire  T_2162_24;
  wire  T_2162_25;
  wire  T_2162_26;
  wire  T_2162_27;
  wire  T_2162_28;
  wire  T_2162_29;
  wire  T_2162_30;
  wire  T_2162_31;
  wire  T_2162_32;
  wire  T_2162_33;
  wire  T_2162_34;
  wire  T_2162_35;
  wire  T_2162_36;
  wire  T_2162_37;
  wire  T_2162_38;
  wire  T_2162_39;
  wire  T_2162_40;
  wire  T_2162_41;
  wire  T_2162_42;
  wire  T_2162_43;
  wire  T_2162_44;
  wire  T_2162_45;
  wire  T_2162_46;
  wire  T_2162_47;
  wire  T_2162_48;
  wire  T_2162_49;
  wire  T_2162_50;
  wire  T_2162_51;
  wire  T_2162_52;
  wire  T_2162_53;
  wire  T_2162_54;
  wire  T_2162_55;
  wire  T_2162_56;
  wire  T_2162_57;
  wire  T_2162_58;
  wire  T_2162_59;
  wire  T_2162_60;
  wire  T_2162_61;
  wire [5:0] T_2225;
  wire [5:0] T_2226;
  wire [5:0] T_2227;
  wire [5:0] T_2228;
  wire [5:0] T_2229;
  wire [5:0] T_2230;
  wire [5:0] T_2231;
  wire [5:0] T_2232;
  wire [5:0] T_2233;
  wire [5:0] T_2234;
  wire [5:0] T_2235;
  wire [5:0] T_2236;
  wire [5:0] T_2237;
  wire [5:0] T_2238;
  wire [5:0] T_2239;
  wire [5:0] T_2240;
  wire [5:0] T_2241;
  wire [5:0] T_2242;
  wire [5:0] T_2243;
  wire [5:0] T_2244;
  wire [5:0] T_2245;
  wire [5:0] T_2246;
  wire [5:0] T_2247;
  wire [5:0] T_2248;
  wire [5:0] T_2249;
  wire [5:0] T_2250;
  wire [5:0] T_2251;
  wire [5:0] T_2252;
  wire [5:0] T_2253;
  wire [5:0] T_2254;
  wire [5:0] T_2255;
  wire [5:0] T_2256;
  wire [5:0] T_2257;
  wire [5:0] T_2258;
  wire [5:0] T_2259;
  wire [5:0] T_2260;
  wire [5:0] T_2261;
  wire [5:0] T_2262;
  wire [5:0] T_2263;
  wire [5:0] T_2264;
  wire [5:0] T_2265;
  wire [5:0] T_2266;
  wire [5:0] T_2267;
  wire [5:0] T_2268;
  wire [5:0] T_2269;
  wire [5:0] T_2270;
  wire [5:0] T_2271;
  wire [5:0] T_2272;
  wire [5:0] T_2273;
  wire [5:0] T_2274;
  wire [5:0] T_2275;
  wire [5:0] T_2276;
  wire [5:0] T_2277;
  wire [5:0] T_2278;
  wire [5:0] T_2279;
  wire [5:0] T_2280;
  wire [5:0] T_2281;
  wire [5:0] T_2282;
  wire [5:0] T_2283;
  wire [5:0] T_2284;
  wire [5:0] T_2285;
  wire [5:0] T_2286;
  wire  T_2288;
  wire  T_2290;
  wire  T_2292;
  wire  T_2294;
  wire  T_2296;
  wire  T_2298;
  wire  T_2300;
  wire  T_2302;
  wire  T_2304;
  wire  T_2306;
  wire  T_2308;
  wire  T_2310;
  wire  T_2312;
  wire  T_2314;
  wire  T_2316;
  wire  T_2318;
  wire  T_2320;
  wire  T_2322;
  wire  T_2324;
  wire  T_2326;
  wire  T_2328;
  wire  T_2330;
  wire  T_2332;
  wire  T_2334;
  wire  T_2336;
  wire  T_2338;
  wire  T_2340;
  wire  T_2342;
  wire  T_2344;
  wire  T_2346;
  wire  T_2348;
  wire  T_2350;
  wire  T_2352;
  wire  T_2354;
  wire  T_2356;
  wire  T_2358;
  wire  T_2360;
  wire  T_2362;
  wire  T_2364;
  wire  T_2366;
  wire  T_2368;
  wire  T_2370;
  wire  T_2372;
  wire  T_2374;
  wire  T_2376;
  wire  T_2378;
  wire  T_2380;
  wire  T_2382;
  wire  T_2384;
  wire  T_2386;
  wire  T_2388;
  wire  T_2390;
  wire  T_2392;
  wire  T_2394;
  wire  T_2396;
  wire  T_2398;
  wire  T_2400;
  wire  T_2402;
  wire  T_2404;
  wire  T_2406;
  wire  T_2408;
  wire  T_2410;
  wire  T_2416_0;
  wire  T_2416_1;
  wire  T_2416_2;
  wire  T_2416_3;
  wire  T_2416_4;
  wire  T_2416_5;
  wire  T_2416_6;
  wire  T_2416_7;
  wire  T_2416_8;
  wire  T_2416_9;
  wire  T_2416_10;
  wire  T_2416_11;
  wire  T_2416_12;
  wire  T_2416_13;
  wire  T_2416_14;
  wire  T_2416_15;
  wire  T_2416_16;
  wire  T_2416_17;
  wire  T_2416_18;
  wire  T_2416_19;
  wire  T_2416_20;
  wire  T_2416_21;
  wire  T_2416_22;
  wire  T_2416_23;
  wire  T_2416_24;
  wire  T_2416_25;
  wire  T_2416_26;
  wire  T_2416_27;
  wire  T_2416_28;
  wire  T_2416_29;
  wire  T_2416_30;
  wire  T_2416_31;
  wire  T_2416_32;
  wire  T_2416_33;
  wire  T_2416_34;
  wire  T_2416_35;
  wire  T_2416_36;
  wire  T_2416_37;
  wire  T_2416_38;
  wire  T_2416_39;
  wire  T_2416_40;
  wire  T_2416_41;
  wire  T_2416_42;
  wire  T_2416_43;
  wire  T_2416_44;
  wire  T_2416_45;
  wire  T_2416_46;
  wire  T_2416_47;
  wire  T_2416_48;
  wire  T_2416_49;
  wire  T_2416_50;
  wire  T_2416_51;
  wire  T_2416_52;
  wire  T_2416_53;
  wire  T_2416_54;
  wire  T_2416_55;
  wire  T_2416_56;
  wire  T_2416_57;
  wire  T_2416_58;
  wire  T_2416_59;
  wire  T_2416_60;
  wire  T_2416_61;
  wire  T_2481;
  wire  T_2482;
  reg [5:0] nextRepl;
  reg [31:0] GEN_430;
  wire  T_2485;
  wire [5:0] GEN_705;
  wire [6:0] T_2487;
  wire [5:0] T_2488;
  wire [5:0] GEN_18;
  wire [5:0] GEN_19;
  wire  useUpdatePageHit;
  wire  doIdxPageRepl;
  wire [5:0] idxPageRepl;
  wire [5:0] idxPageUpdateOH;
  wire [1:0] T_2494;
  wire [3:0] T_2495;
  wire [1:0] GEN_707;
  wire  T_2497;
  wire [3:0] GEN_708;
  wire [3:0] T_2498;
  wire [1:0] T_2499;
  wire [1:0] T_2500;
  wire  T_2502;
  wire [1:0] T_2503;
  wire  T_2504;
  wire [1:0] T_2505;
  wire [2:0] idxPageUpdate;
  wire [5:0] idxPageReplEn;
  wire  samePage;
  wire [5:0] T_2509;
  wire [5:0] T_2510;
  wire  usePageHit;
  wire  T_2513;
  wire  T_2515;
  wire  doTgtPageRepl;
  wire [4:0] T_2516;
  wire [5:0] GEN_711;
  wire [5:0] T_2517;
  wire  T_2518;
  wire [5:0] GEN_712;
  wire [5:0] T_2519;
  wire [5:0] tgtPageRepl;
  wire [5:0] T_2520;
  wire [1:0] T_2521;
  wire [3:0] T_2522;
  wire  T_2524;
  wire [3:0] GEN_714;
  wire [3:0] T_2525;
  wire [1:0] T_2526;
  wire [1:0] T_2527;
  wire  T_2529;
  wire [1:0] T_2530;
  wire  T_2531;
  wire [1:0] T_2532;
  wire [2:0] tgtPageUpdate;
  wire [5:0] tgtPageReplEn;
  wire  doPageRepl;
  wire [5:0] pageReplEn;
  wire  T_2534;
  reg [2:0] T_2536;
  reg [31:0] GEN_434;
  wire  T_2538;
  wire [2:0] GEN_716;
  wire [3:0] T_2540;
  wire [2:0] T_2541;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire [7:0] T_2545;
  wire  T_2546;
  wire  T_2547;
  wire  T_2549;
  wire [5:0] T_2550;
  wire [5:0] T_2551;
  wire [5:0] T_2552;
  wire  T_2554;
  wire [5:0] T_2555;
  wire [5:0] T_2556;
  wire  T_2558;
  wire [5:0] T_2559;
  wire [5:0] T_2560;
  wire  T_2562;
  wire [5:0] T_2563;
  wire [5:0] T_2564;
  wire  T_2566;
  wire [5:0] T_2567;
  wire [5:0] T_2568;
  wire  T_2570;
  wire [5:0] T_2571;
  wire [5:0] T_2572;
  wire  T_2574;
  wire [5:0] T_2575;
  wire [5:0] T_2576;
  wire  T_2578;
  wire [5:0] T_2579;
  wire [5:0] T_2580;
  wire  T_2582;
  wire [5:0] T_2583;
  wire [5:0] T_2584;
  wire  T_2586;
  wire [5:0] T_2587;
  wire [5:0] T_2588;
  wire  T_2590;
  wire [5:0] T_2591;
  wire [5:0] T_2592;
  wire  T_2594;
  wire [5:0] T_2595;
  wire [5:0] T_2596;
  wire  T_2598;
  wire [5:0] T_2599;
  wire [5:0] T_2600;
  wire  T_2602;
  wire [5:0] T_2603;
  wire [5:0] T_2604;
  wire  T_2606;
  wire [5:0] T_2607;
  wire [5:0] T_2608;
  wire  T_2610;
  wire [5:0] T_2611;
  wire [5:0] T_2612;
  wire  T_2614;
  wire [5:0] T_2615;
  wire [5:0] T_2616;
  wire  T_2618;
  wire [5:0] T_2619;
  wire [5:0] T_2620;
  wire  T_2622;
  wire [5:0] T_2623;
  wire [5:0] T_2624;
  wire  T_2626;
  wire [5:0] T_2627;
  wire [5:0] T_2628;
  wire  T_2630;
  wire [5:0] T_2631;
  wire [5:0] T_2632;
  wire  T_2634;
  wire [5:0] T_2635;
  wire [5:0] T_2636;
  wire  T_2638;
  wire [5:0] T_2639;
  wire [5:0] T_2640;
  wire  T_2642;
  wire [5:0] T_2643;
  wire [5:0] T_2644;
  wire  T_2646;
  wire [5:0] T_2647;
  wire [5:0] T_2648;
  wire  T_2650;
  wire [5:0] T_2651;
  wire [5:0] T_2652;
  wire  T_2654;
  wire [5:0] T_2655;
  wire [5:0] T_2656;
  wire  T_2658;
  wire [5:0] T_2659;
  wire [5:0] T_2660;
  wire  T_2662;
  wire [5:0] T_2663;
  wire [5:0] T_2664;
  wire  T_2666;
  wire [5:0] T_2667;
  wire [5:0] T_2668;
  wire  T_2670;
  wire [5:0] T_2671;
  wire [5:0] T_2672;
  wire  T_2674;
  wire [5:0] T_2675;
  wire [5:0] T_2676;
  wire  T_2678;
  wire [5:0] T_2679;
  wire [5:0] T_2680;
  wire  T_2682;
  wire [5:0] T_2683;
  wire [5:0] T_2684;
  wire  T_2686;
  wire [5:0] T_2687;
  wire [5:0] T_2688;
  wire  T_2690;
  wire [5:0] T_2691;
  wire [5:0] T_2692;
  wire  T_2694;
  wire [5:0] T_2695;
  wire [5:0] T_2696;
  wire  T_2698;
  wire [5:0] T_2699;
  wire [5:0] T_2700;
  wire  T_2702;
  wire [5:0] T_2703;
  wire [5:0] T_2704;
  wire  T_2706;
  wire [5:0] T_2707;
  wire [5:0] T_2708;
  wire  T_2710;
  wire [5:0] T_2711;
  wire [5:0] T_2712;
  wire  T_2714;
  wire [5:0] T_2715;
  wire [5:0] T_2716;
  wire  T_2718;
  wire [5:0] T_2719;
  wire [5:0] T_2720;
  wire  T_2722;
  wire [5:0] T_2723;
  wire [5:0] T_2724;
  wire  T_2726;
  wire [5:0] T_2727;
  wire [5:0] T_2728;
  wire  T_2730;
  wire [5:0] T_2731;
  wire [5:0] T_2732;
  wire  T_2734;
  wire [5:0] T_2735;
  wire [5:0] T_2736;
  wire  T_2738;
  wire [5:0] T_2739;
  wire [5:0] T_2740;
  wire  T_2742;
  wire [5:0] T_2743;
  wire [5:0] T_2744;
  wire  T_2746;
  wire [5:0] T_2747;
  wire [5:0] T_2748;
  wire  T_2750;
  wire [5:0] T_2751;
  wire [5:0] T_2752;
  wire  T_2754;
  wire [5:0] T_2755;
  wire [5:0] T_2756;
  wire  T_2758;
  wire [5:0] T_2759;
  wire [5:0] T_2760;
  wire  T_2762;
  wire [5:0] T_2763;
  wire [5:0] T_2764;
  wire  T_2766;
  wire [5:0] T_2767;
  wire [5:0] T_2768;
  wire  T_2770;
  wire [5:0] T_2771;
  wire [5:0] T_2772;
  wire  T_2774;
  wire [5:0] T_2775;
  wire [5:0] T_2776;
  wire  T_2778;
  wire [5:0] T_2779;
  wire [5:0] T_2780;
  wire  T_2782;
  wire [5:0] T_2783;
  wire [5:0] T_2784;
  wire  T_2786;
  wire [5:0] T_2787;
  wire [5:0] T_2788;
  wire  T_2790;
  wire [5:0] T_2791;
  wire [5:0] T_2792;
  wire  T_2794;
  wire [5:0] T_2795;
  wire [5:0] T_2796;
  wire  T_2798;
  wire  T_2804_0;
  wire  T_2804_1;
  wire  T_2804_2;
  wire  T_2804_3;
  wire  T_2804_4;
  wire  T_2804_5;
  wire  T_2804_6;
  wire  T_2804_7;
  wire  T_2804_8;
  wire  T_2804_9;
  wire  T_2804_10;
  wire  T_2804_11;
  wire  T_2804_12;
  wire  T_2804_13;
  wire  T_2804_14;
  wire  T_2804_15;
  wire  T_2804_16;
  wire  T_2804_17;
  wire  T_2804_18;
  wire  T_2804_19;
  wire  T_2804_20;
  wire  T_2804_21;
  wire  T_2804_22;
  wire  T_2804_23;
  wire  T_2804_24;
  wire  T_2804_25;
  wire  T_2804_26;
  wire  T_2804_27;
  wire  T_2804_28;
  wire  T_2804_29;
  wire  T_2804_30;
  wire  T_2804_31;
  wire  T_2804_32;
  wire  T_2804_33;
  wire  T_2804_34;
  wire  T_2804_35;
  wire  T_2804_36;
  wire  T_2804_37;
  wire  T_2804_38;
  wire  T_2804_39;
  wire  T_2804_40;
  wire  T_2804_41;
  wire  T_2804_42;
  wire  T_2804_43;
  wire  T_2804_44;
  wire  T_2804_45;
  wire  T_2804_46;
  wire  T_2804_47;
  wire  T_2804_48;
  wire  T_2804_49;
  wire  T_2804_50;
  wire  T_2804_51;
  wire  T_2804_52;
  wire  T_2804_53;
  wire  T_2804_54;
  wire  T_2804_55;
  wire  T_2804_56;
  wire  T_2804_57;
  wire  T_2804_58;
  wire  T_2804_59;
  wire  T_2804_60;
  wire  T_2804_61;
  wire [1:0] T_2806;
  wire [2:0] T_2807;
  wire [1:0] T_2808;
  wire [1:0] T_2809;
  wire [3:0] T_2810;
  wire [6:0] T_2811;
  wire [1:0] T_2812;
  wire [1:0] T_2813;
  wire [3:0] T_2814;
  wire [1:0] T_2815;
  wire [1:0] T_2816;
  wire [3:0] T_2817;
  wire [7:0] T_2818;
  wire [14:0] T_2819;
  wire [1:0] T_2820;
  wire [1:0] T_2821;
  wire [3:0] T_2822;
  wire [1:0] T_2823;
  wire [1:0] T_2824;
  wire [3:0] T_2825;
  wire [7:0] T_2826;
  wire [1:0] T_2827;
  wire [1:0] T_2828;
  wire [3:0] T_2829;
  wire [1:0] T_2830;
  wire [1:0] T_2831;
  wire [3:0] T_2832;
  wire [7:0] T_2833;
  wire [15:0] T_2834;
  wire [30:0] T_2835;
  wire [1:0] T_2836;
  wire [2:0] T_2837;
  wire [1:0] T_2838;
  wire [1:0] T_2839;
  wire [3:0] T_2840;
  wire [6:0] T_2841;
  wire [1:0] T_2842;
  wire [1:0] T_2843;
  wire [3:0] T_2844;
  wire [1:0] T_2845;
  wire [1:0] T_2846;
  wire [3:0] T_2847;
  wire [7:0] T_2848;
  wire [14:0] T_2849;
  wire [1:0] T_2850;
  wire [1:0] T_2851;
  wire [3:0] T_2852;
  wire [1:0] T_2853;
  wire [1:0] T_2854;
  wire [3:0] T_2855;
  wire [7:0] T_2856;
  wire [1:0] T_2857;
  wire [1:0] T_2858;
  wire [3:0] T_2859;
  wire [1:0] T_2860;
  wire [1:0] T_2861;
  wire [3:0] T_2862;
  wire [7:0] T_2863;
  wire [15:0] T_2864;
  wire [30:0] T_2865;
  wire [61:0] T_2866;
  wire [63:0] GEN_780;
  wire [63:0] T_2868;
  wire [61:0] T_2869;
  wire [61:0] T_2870;
  wire [63:0] GEN_781;
  wire [63:0] T_2871;
  wire  GEN_0;
  wire  GEN_22;
  wire  GEN_23;
  wire [5:0] GEN_784;
  wire  GEN_24;
  wire [5:0] GEN_785;
  wire  GEN_25;
  wire [5:0] GEN_786;
  wire  GEN_26;
  wire [5:0] GEN_787;
  wire  GEN_27;
  wire [5:0] GEN_788;
  wire  GEN_28;
  wire [5:0] GEN_789;
  wire  GEN_29;
  wire [5:0] GEN_790;
  wire  GEN_30;
  wire [5:0] GEN_791;
  wire  GEN_31;
  wire [5:0] GEN_792;
  wire  GEN_32;
  wire [5:0] GEN_793;
  wire  GEN_33;
  wire [5:0] GEN_794;
  wire  GEN_34;
  wire [5:0] GEN_795;
  wire  GEN_35;
  wire [5:0] GEN_796;
  wire  GEN_36;
  wire [5:0] GEN_797;
  wire  GEN_37;
  wire [5:0] GEN_798;
  wire  GEN_38;
  wire [5:0] GEN_799;
  wire  GEN_39;
  wire [5:0] GEN_800;
  wire  GEN_40;
  wire [5:0] GEN_801;
  wire  GEN_41;
  wire [5:0] GEN_802;
  wire  GEN_42;
  wire [5:0] GEN_803;
  wire  GEN_43;
  wire [5:0] GEN_804;
  wire  GEN_44;
  wire [5:0] GEN_805;
  wire  GEN_45;
  wire [5:0] GEN_806;
  wire  GEN_46;
  wire [5:0] GEN_807;
  wire  GEN_47;
  wire [5:0] GEN_808;
  wire  GEN_48;
  wire [5:0] GEN_809;
  wire  GEN_49;
  wire [5:0] GEN_810;
  wire  GEN_50;
  wire [5:0] GEN_811;
  wire  GEN_51;
  wire [5:0] GEN_812;
  wire  GEN_52;
  wire [5:0] GEN_813;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire  GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_62;
  wire  GEN_63;
  wire  GEN_64;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_1;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire [5:0] T_2881;
  wire  T_2883;
  wire  T_2884;
  wire [26:0] T_2887;
  wire  T_2888;
  wire  T_2889;
  wire  T_2892;
  wire  T_2893;
  wire  T_2896;
  wire  T_2897;
  wire  T_2900;
  wire [26:0] T_2903;
  wire  T_2904;
  wire  T_2905;
  wire  T_2908;
  wire  T_2909;
  wire  T_2912;
  wire  T_2913;
  wire [5:0] T_2916;
  wire [5:0] GEN_176;
  wire [63:0] GEN_239;
  wire  GEN_261;
  wire  GEN_262;
  wire  GEN_263;
  wire  GEN_264;
  wire  GEN_265;
  wire  GEN_266;
  wire  GEN_267;
  wire  GEN_268;
  wire  GEN_269;
  wire  GEN_270;
  wire  GEN_271;
  wire  GEN_272;
  wire  GEN_273;
  wire  GEN_274;
  wire  GEN_275;
  wire  GEN_276;
  wire  GEN_277;
  wire  GEN_278;
  wire  GEN_279;
  wire  GEN_280;
  wire  GEN_281;
  wire  GEN_282;
  wire  GEN_283;
  wire  GEN_284;
  wire  GEN_285;
  wire  GEN_286;
  wire  GEN_287;
  wire  GEN_288;
  wire  GEN_289;
  wire  GEN_290;
  wire  GEN_291;
  wire  GEN_292;
  wire  GEN_293;
  wire  GEN_294;
  wire  GEN_295;
  wire  GEN_296;
  wire  GEN_297;
  wire  GEN_298;
  wire  GEN_299;
  wire  GEN_300;
  wire  GEN_301;
  wire  GEN_302;
  wire  GEN_303;
  wire  GEN_304;
  wire  GEN_305;
  wire  GEN_306;
  wire  GEN_307;
  wire  GEN_308;
  wire  GEN_309;
  wire  GEN_310;
  wire  GEN_311;
  wire  GEN_312;
  wire  GEN_313;
  wire  GEN_314;
  wire  GEN_315;
  wire  GEN_316;
  wire  GEN_317;
  wire  GEN_318;
  wire  GEN_319;
  wire  GEN_320;
  wire  GEN_321;
  wire  GEN_322;
  wire  GEN_324;
  wire  GEN_325;
  wire  GEN_326;
  wire  GEN_327;
  wire  GEN_328;
  wire  GEN_329;
  wire  GEN_330;
  wire  GEN_331;
  wire  GEN_332;
  wire  GEN_333;
  wire  GEN_334;
  wire  GEN_335;
  wire  GEN_336;
  wire  GEN_337;
  wire  GEN_338;
  wire  GEN_339;
  wire  GEN_340;
  wire  GEN_341;
  wire  GEN_342;
  wire  GEN_343;
  wire  GEN_344;
  wire  GEN_345;
  wire  GEN_346;
  wire  GEN_347;
  wire  GEN_348;
  wire  GEN_349;
  wire  GEN_350;
  wire  GEN_351;
  wire  GEN_352;
  wire  GEN_353;
  wire  GEN_354;
  wire  GEN_355;
  wire  GEN_356;
  wire  GEN_357;
  wire  GEN_358;
  wire  GEN_359;
  wire  GEN_360;
  wire  GEN_361;
  wire  GEN_362;
  wire  GEN_363;
  wire  GEN_364;
  wire  GEN_365;
  wire  GEN_366;
  wire  GEN_367;
  wire  GEN_368;
  wire  GEN_369;
  wire  GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire  GEN_373;
  wire  GEN_374;
  wire  GEN_375;
  wire  GEN_376;
  wire  GEN_377;
  wire  GEN_378;
  wire  GEN_379;
  wire  GEN_380;
  wire  GEN_381;
  wire  GEN_382;
  wire  GEN_383;
  wire  GEN_384;
  wire  GEN_385;
  wire  GEN_393;
  wire  GEN_398;
  wire  GEN_403;
  wire  GEN_408;
  wire  GEN_413;
  wire  GEN_418;
  wire [5:0] GEN_421;
  wire [63:0] GEN_422;
  wire [5:0] GEN_423;
  wire [61:0] GEN_847;
  wire  T_2920;
  wire  T_2921;
  wire  T_2922;
  wire  T_2923;
  wire  T_2924;
  wire  T_2925;
  wire  T_2926;
  wire  T_2927;
  wire  T_2928;
  wire  T_2929;
  wire  T_2930;
  wire  T_2931;
  wire  T_2932;
  wire  T_2933;
  wire  T_2934;
  wire  T_2935;
  wire  T_2936;
  wire  T_2937;
  wire  T_2938;
  wire  T_2939;
  wire  T_2940;
  wire  T_2941;
  wire  T_2942;
  wire  T_2943;
  wire  T_2944;
  wire  T_2945;
  wire  T_2946;
  wire  T_2947;
  wire  T_2948;
  wire  T_2949;
  wire  T_2950;
  wire  T_2951;
  wire  T_2952;
  wire  T_2953;
  wire  T_2954;
  wire  T_2955;
  wire  T_2956;
  wire  T_2957;
  wire  T_2958;
  wire  T_2959;
  wire  T_2960;
  wire  T_2961;
  wire  T_2962;
  wire  T_2963;
  wire  T_2964;
  wire  T_2965;
  wire  T_2966;
  wire  T_2967;
  wire  T_2968;
  wire  T_2969;
  wire  T_2970;
  wire  T_2971;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2977;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2981;
  wire  T_2982;
  wire [5:0] T_2984;
  wire [5:0] T_2986;
  wire [5:0] T_2988;
  wire [5:0] T_2990;
  wire [5:0] T_2992;
  wire [5:0] T_2994;
  wire [5:0] T_2996;
  wire [5:0] T_2998;
  wire [5:0] T_3000;
  wire [5:0] T_3002;
  wire [5:0] T_3004;
  wire [5:0] T_3006;
  wire [5:0] T_3008;
  wire [5:0] T_3010;
  wire [5:0] T_3012;
  wire [5:0] T_3014;
  wire [5:0] T_3016;
  wire [5:0] T_3018;
  wire [5:0] T_3020;
  wire [5:0] T_3022;
  wire [5:0] T_3024;
  wire [5:0] T_3026;
  wire [5:0] T_3028;
  wire [5:0] T_3030;
  wire [5:0] T_3032;
  wire [5:0] T_3034;
  wire [5:0] T_3036;
  wire [5:0] T_3038;
  wire [5:0] T_3040;
  wire [5:0] T_3042;
  wire [5:0] T_3044;
  wire [5:0] T_3046;
  wire [5:0] T_3048;
  wire [5:0] T_3050;
  wire [5:0] T_3052;
  wire [5:0] T_3054;
  wire [5:0] T_3056;
  wire [5:0] T_3058;
  wire [5:0] T_3060;
  wire [5:0] T_3062;
  wire [5:0] T_3064;
  wire [5:0] T_3066;
  wire [5:0] T_3068;
  wire [5:0] T_3070;
  wire [5:0] T_3072;
  wire [5:0] T_3074;
  wire [5:0] T_3076;
  wire [5:0] T_3078;
  wire [5:0] T_3080;
  wire [5:0] T_3082;
  wire [5:0] T_3084;
  wire [5:0] T_3086;
  wire [5:0] T_3088;
  wire [5:0] T_3090;
  wire [5:0] T_3092;
  wire [5:0] T_3094;
  wire [5:0] T_3096;
  wire [5:0] T_3098;
  wire [5:0] T_3100;
  wire [5:0] T_3102;
  wire [5:0] T_3104;
  wire [5:0] T_3106;
  wire [5:0] T_3108;
  wire [5:0] T_3109;
  wire [5:0] T_3110;
  wire [5:0] T_3111;
  wire [5:0] T_3112;
  wire [5:0] T_3113;
  wire [5:0] T_3114;
  wire [5:0] T_3115;
  wire [5:0] T_3116;
  wire [5:0] T_3117;
  wire [5:0] T_3118;
  wire [5:0] T_3119;
  wire [5:0] T_3120;
  wire [5:0] T_3121;
  wire [5:0] T_3122;
  wire [5:0] T_3123;
  wire [5:0] T_3124;
  wire [5:0] T_3125;
  wire [5:0] T_3126;
  wire [5:0] T_3127;
  wire [5:0] T_3128;
  wire [5:0] T_3129;
  wire [5:0] T_3130;
  wire [5:0] T_3131;
  wire [5:0] T_3132;
  wire [5:0] T_3133;
  wire [5:0] T_3134;
  wire [5:0] T_3135;
  wire [5:0] T_3136;
  wire [5:0] T_3137;
  wire [5:0] T_3138;
  wire [5:0] T_3139;
  wire [5:0] T_3140;
  wire [5:0] T_3141;
  wire [5:0] T_3142;
  wire [5:0] T_3143;
  wire [5:0] T_3144;
  wire [5:0] T_3145;
  wire [5:0] T_3146;
  wire [5:0] T_3147;
  wire [5:0] T_3148;
  wire [5:0] T_3149;
  wire [5:0] T_3150;
  wire [5:0] T_3151;
  wire [5:0] T_3152;
  wire [5:0] T_3153;
  wire [5:0] T_3154;
  wire [5:0] T_3155;
  wire [5:0] T_3156;
  wire [5:0] T_3157;
  wire [5:0] T_3158;
  wire [5:0] T_3159;
  wire [5:0] T_3160;
  wire [5:0] T_3161;
  wire [5:0] T_3162;
  wire [5:0] T_3163;
  wire [5:0] T_3164;
  wire [5:0] T_3165;
  wire [5:0] T_3166;
  wire [5:0] T_3167;
  wire [5:0] T_3168;
  wire [5:0] T_3169;
  wire  T_3170;
  wire  T_3171;
  wire  T_3172;
  wire  T_3173;
  wire  T_3174;
  wire  T_3175;
  wire [26:0] T_3189;
  wire [26:0] T_3191;
  wire [26:0] T_3193;
  wire [26:0] T_3195;
  wire [26:0] T_3197;
  wire [26:0] T_3199;
  wire [26:0] T_3201;
  wire [26:0] T_3202;
  wire [26:0] T_3203;
  wire [26:0] T_3204;
  wire [26:0] T_3205;
  wire [26:0] T_3206;
  wire [11:0] T_3394;
  wire [11:0] T_3396;
  wire [11:0] T_3398;
  wire [11:0] T_3400;
  wire [11:0] T_3402;
  wire [11:0] T_3404;
  wire [11:0] T_3406;
  wire [11:0] T_3408;
  wire [11:0] T_3410;
  wire [11:0] T_3412;
  wire [11:0] T_3414;
  wire [11:0] T_3416;
  wire [11:0] T_3418;
  wire [11:0] T_3420;
  wire [11:0] T_3422;
  wire [11:0] T_3424;
  wire [11:0] T_3426;
  wire [11:0] T_3428;
  wire [11:0] T_3430;
  wire [11:0] T_3432;
  wire [11:0] T_3434;
  wire [11:0] T_3436;
  wire [11:0] T_3438;
  wire [11:0] T_3440;
  wire [11:0] T_3442;
  wire [11:0] T_3444;
  wire [11:0] T_3446;
  wire [11:0] T_3448;
  wire [11:0] T_3450;
  wire [11:0] T_3452;
  wire [11:0] T_3454;
  wire [11:0] T_3456;
  wire [11:0] T_3458;
  wire [11:0] T_3460;
  wire [11:0] T_3462;
  wire [11:0] T_3464;
  wire [11:0] T_3466;
  wire [11:0] T_3468;
  wire [11:0] T_3470;
  wire [11:0] T_3472;
  wire [11:0] T_3474;
  wire [11:0] T_3476;
  wire [11:0] T_3478;
  wire [11:0] T_3480;
  wire [11:0] T_3482;
  wire [11:0] T_3484;
  wire [11:0] T_3486;
  wire [11:0] T_3488;
  wire [11:0] T_3490;
  wire [11:0] T_3492;
  wire [11:0] T_3494;
  wire [11:0] T_3496;
  wire [11:0] T_3498;
  wire [11:0] T_3500;
  wire [11:0] T_3502;
  wire [11:0] T_3504;
  wire [11:0] T_3506;
  wire [11:0] T_3508;
  wire [11:0] T_3510;
  wire [11:0] T_3512;
  wire [11:0] T_3514;
  wire [11:0] T_3516;
  wire [11:0] T_3518;
  wire [11:0] T_3519;
  wire [11:0] T_3520;
  wire [11:0] T_3521;
  wire [11:0] T_3522;
  wire [11:0] T_3523;
  wire [11:0] T_3524;
  wire [11:0] T_3525;
  wire [11:0] T_3526;
  wire [11:0] T_3527;
  wire [11:0] T_3528;
  wire [11:0] T_3529;
  wire [11:0] T_3530;
  wire [11:0] T_3531;
  wire [11:0] T_3532;
  wire [11:0] T_3533;
  wire [11:0] T_3534;
  wire [11:0] T_3535;
  wire [11:0] T_3536;
  wire [11:0] T_3537;
  wire [11:0] T_3538;
  wire [11:0] T_3539;
  wire [11:0] T_3540;
  wire [11:0] T_3541;
  wire [11:0] T_3542;
  wire [11:0] T_3543;
  wire [11:0] T_3544;
  wire [11:0] T_3545;
  wire [11:0] T_3546;
  wire [11:0] T_3547;
  wire [11:0] T_3548;
  wire [11:0] T_3549;
  wire [11:0] T_3550;
  wire [11:0] T_3551;
  wire [11:0] T_3552;
  wire [11:0] T_3553;
  wire [11:0] T_3554;
  wire [11:0] T_3555;
  wire [11:0] T_3556;
  wire [11:0] T_3557;
  wire [11:0] T_3558;
  wire [11:0] T_3559;
  wire [11:0] T_3560;
  wire [11:0] T_3561;
  wire [11:0] T_3562;
  wire [11:0] T_3563;
  wire [11:0] T_3564;
  wire [11:0] T_3565;
  wire [11:0] T_3566;
  wire [11:0] T_3567;
  wire [11:0] T_3568;
  wire [11:0] T_3569;
  wire [11:0] T_3570;
  wire [11:0] T_3571;
  wire [11:0] T_3572;
  wire [11:0] T_3573;
  wire [11:0] T_3574;
  wire [11:0] T_3575;
  wire [11:0] T_3576;
  wire [11:0] T_3577;
  wire [11:0] T_3578;
  wire [11:0] T_3579;
  wire [38:0] T_3580;
  wire [29:0] T_3581;
  wire [31:0] T_3582;
  wire [29:0] GEN_848;
  wire  T_3584;
  wire [31:0] GEN_849;
  wire [31:0] T_3585;
  wire [15:0] T_3586;
  wire [15:0] T_3587;
  wire [15:0] GEN_850;
  wire  T_3589;
  wire [15:0] T_3590;
  wire [7:0] T_3591;
  wire [7:0] T_3592;
  wire [7:0] GEN_851;
  wire  T_3594;
  wire [7:0] T_3595;
  wire [3:0] T_3596;
  wire [3:0] T_3597;
  wire [3:0] GEN_852;
  wire  T_3599;
  wire [3:0] T_3600;
  wire [1:0] T_3601;
  wire [1:0] T_3602;
  wire  T_3604;
  wire [1:0] T_3605;
  wire  T_3606;
  wire [1:0] T_3607;
  wire [2:0] T_3608;
  wire [3:0] T_3609;
  wire [4:0] T_3610;
  wire [5:0] T_3611;
  reg [1:0] T_3616 [0:127];
  reg [31:0] GEN_441;
  wire [1:0] T_3616_T_3942_data;
  wire [6:0] T_3616_T_3942_addr;
  wire  T_3616_T_3942_en;
  wire [1:0] T_3616_T_3949_data;
  wire [6:0] T_3616_T_3949_addr;
  wire  T_3616_T_3949_mask;
  wire  T_3616_T_3949_en;
  reg [6:0] T_3618;
  reg [31:0] GEN_451;
  wire  T_3683;
  wire  T_3686;
  wire  T_3689;
  wire  T_3692;
  wire  T_3695;
  wire  T_3698;
  wire  T_3701;
  wire  T_3704;
  wire  T_3707;
  wire  T_3710;
  wire  T_3713;
  wire  T_3716;
  wire  T_3719;
  wire  T_3722;
  wire  T_3725;
  wire  T_3728;
  wire  T_3731;
  wire  T_3734;
  wire  T_3737;
  wire  T_3740;
  wire  T_3743;
  wire  T_3746;
  wire  T_3749;
  wire  T_3752;
  wire  T_3755;
  wire  T_3758;
  wire  T_3761;
  wire  T_3764;
  wire  T_3767;
  wire  T_3770;
  wire  T_3773;
  wire  T_3776;
  wire  T_3779;
  wire  T_3782;
  wire  T_3785;
  wire  T_3788;
  wire  T_3791;
  wire  T_3794;
  wire  T_3797;
  wire  T_3800;
  wire  T_3803;
  wire  T_3806;
  wire  T_3809;
  wire  T_3812;
  wire  T_3815;
  wire  T_3818;
  wire  T_3821;
  wire  T_3824;
  wire  T_3827;
  wire  T_3830;
  wire  T_3833;
  wire  T_3836;
  wire  T_3839;
  wire  T_3842;
  wire  T_3845;
  wire  T_3848;
  wire  T_3851;
  wire  T_3854;
  wire  T_3857;
  wire  T_3860;
  wire  T_3863;
  wire  T_3866;
  wire  T_3868;
  wire  T_3869;
  wire  T_3870;
  wire  T_3871;
  wire  T_3872;
  wire  T_3873;
  wire  T_3874;
  wire  T_3875;
  wire  T_3876;
  wire  T_3877;
  wire  T_3878;
  wire  T_3879;
  wire  T_3880;
  wire  T_3881;
  wire  T_3882;
  wire  T_3883;
  wire  T_3884;
  wire  T_3885;
  wire  T_3886;
  wire  T_3887;
  wire  T_3888;
  wire  T_3889;
  wire  T_3890;
  wire  T_3891;
  wire  T_3892;
  wire  T_3893;
  wire  T_3894;
  wire  T_3895;
  wire  T_3896;
  wire  T_3897;
  wire  T_3898;
  wire  T_3899;
  wire  T_3900;
  wire  T_3901;
  wire  T_3902;
  wire  T_3903;
  wire  T_3904;
  wire  T_3905;
  wire  T_3906;
  wire  T_3907;
  wire  T_3908;
  wire  T_3909;
  wire  T_3910;
  wire  T_3911;
  wire  T_3912;
  wire  T_3913;
  wire  T_3914;
  wire  T_3915;
  wire  T_3916;
  wire  T_3917;
  wire  T_3918;
  wire  T_3919;
  wire  T_3920;
  wire  T_3921;
  wire  T_3922;
  wire  T_3923;
  wire  T_3924;
  wire  T_3925;
  wire  T_3926;
  wire  T_3927;
  wire  T_3928;
  wire  T_3929;
  wire  T_3931;
  wire  T_3932;
  wire  T_3933;
  wire [6:0] T_3937_history;
  wire [1:0] T_3937_value;
  wire [6:0] T_3940;
  wire [6:0] T_3941;
  wire  T_3943;
  wire [5:0] T_3944;
  wire [6:0] T_3945;
  wire [6:0] GEN_424;
  wire  T_3946;
  wire [6:0] T_3947;
  wire [6:0] T_3948;
  wire  T_3950;
  wire  T_3951;
  wire  T_3952;
  wire  T_3955;
  wire  T_3956;
  wire  T_3957;
  wire [1:0] T_3958;
  wire [5:0] T_3959;
  wire [6:0] T_3960;
  wire [6:0] GEN_425;
  wire [6:0] GEN_431;
  wire  T_3963;
  wire  T_3964;
  wire  GEN_432;
  reg [1:0] T_3967;
  reg [31:0] GEN_458;
  reg  T_3969;
  reg [31:0] GEN_459;
  reg [38:0] T_3976_0;
  reg [63:0] GEN_460;
  reg [38:0] T_3976_1;
  reg [63:0] GEN_461;
  wire  T_4042;
  wire  T_4045;
  wire  T_4048;
  wire  T_4051;
  wire  T_4054;
  wire  T_4057;
  wire  T_4060;
  wire  T_4063;
  wire  T_4066;
  wire  T_4069;
  wire  T_4072;
  wire  T_4075;
  wire  T_4078;
  wire  T_4081;
  wire  T_4084;
  wire  T_4087;
  wire  T_4090;
  wire  T_4093;
  wire  T_4096;
  wire  T_4099;
  wire  T_4102;
  wire  T_4105;
  wire  T_4108;
  wire  T_4111;
  wire  T_4114;
  wire  T_4117;
  wire  T_4120;
  wire  T_4123;
  wire  T_4126;
  wire  T_4129;
  wire  T_4132;
  wire  T_4135;
  wire  T_4138;
  wire  T_4141;
  wire  T_4144;
  wire  T_4147;
  wire  T_4150;
  wire  T_4153;
  wire  T_4156;
  wire  T_4159;
  wire  T_4162;
  wire  T_4165;
  wire  T_4168;
  wire  T_4171;
  wire  T_4174;
  wire  T_4177;
  wire  T_4180;
  wire  T_4183;
  wire  T_4186;
  wire  T_4189;
  wire  T_4192;
  wire  T_4195;
  wire  T_4198;
  wire  T_4201;
  wire  T_4204;
  wire  T_4207;
  wire  T_4210;
  wire  T_4213;
  wire  T_4216;
  wire  T_4219;
  wire  T_4222;
  wire  T_4225;
  wire  T_4227;
  wire  T_4228;
  wire  T_4229;
  wire  T_4230;
  wire  T_4231;
  wire  T_4232;
  wire  T_4233;
  wire  T_4234;
  wire  T_4235;
  wire  T_4236;
  wire  T_4237;
  wire  T_4238;
  wire  T_4239;
  wire  T_4240;
  wire  T_4241;
  wire  T_4242;
  wire  T_4243;
  wire  T_4244;
  wire  T_4245;
  wire  T_4246;
  wire  T_4247;
  wire  T_4248;
  wire  T_4249;
  wire  T_4250;
  wire  T_4251;
  wire  T_4252;
  wire  T_4253;
  wire  T_4254;
  wire  T_4255;
  wire  T_4256;
  wire  T_4257;
  wire  T_4258;
  wire  T_4259;
  wire  T_4260;
  wire  T_4261;
  wire  T_4262;
  wire  T_4263;
  wire  T_4264;
  wire  T_4265;
  wire  T_4266;
  wire  T_4267;
  wire  T_4268;
  wire  T_4269;
  wire  T_4270;
  wire  T_4271;
  wire  T_4272;
  wire  T_4273;
  wire  T_4274;
  wire  T_4275;
  wire  T_4276;
  wire  T_4277;
  wire  T_4278;
  wire  T_4279;
  wire  T_4280;
  wire  T_4281;
  wire  T_4282;
  wire  T_4283;
  wire  T_4284;
  wire  T_4285;
  wire  T_4286;
  wire  T_4287;
  wire  T_4288;
  wire  T_4290;
  wire  T_4292;
  wire  T_4293;
  wire [38:0] GEN_2;
  wire [38:0] GEN_433;
  wire [38:0] GEN_435;
  wire  T_4295;
  wire [1:0] GEN_855;
  wire [2:0] T_4297;
  wire [1:0] T_4298;
  wire [1:0] GEN_436;
  wire [1:0] T_4304;
  wire  T_4305;
  wire [38:0] GEN_3;
  wire [38:0] GEN_437;
  wire [38:0] GEN_438;
  wire [38:0] GEN_439;
  wire [1:0] GEN_440;
  wire [38:0] GEN_442;
  wire [38:0] GEN_443;
  wire  GEN_444;
  wire [38:0] GEN_445;
  wire  T_4308;
  wire  T_4310;
  wire  T_4311;
  wire [2:0] T_4317;
  wire [1:0] T_4318;
  wire [1:0] T_4324;
  wire  T_4325;
  wire [1:0] GEN_446;
  wire  GEN_447;
  wire [1:0] GEN_448;
  wire  GEN_449;
  wire [1:0] GEN_450;
  wire [38:0] GEN_452;
  wire [38:0] GEN_453;
  wire  GEN_454;
  wire [38:0] GEN_455;
  wire [1:0] GEN_456;
  assign io_resp_valid = T_2920;
  assign io_resp_bits_taken = GEN_432;
  assign io_resp_bits_mask = 1'h1;
  assign io_resp_bits_bridx = brIdx_T_3612_data;
  assign io_resp_bits_target = GEN_455;
  assign io_resp_bits_entry = T_3611;
  assign io_resp_bits_bht_history = T_3937_history;
  assign io_resp_bits_bht_value = T_3937_value;
  assign idxs_T_1431_addr = {{5'd0}, 1'h0};
  assign idxs_T_1431_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1431_data = idxs[idxs_T_1431_addr];
  `else
  assign idxs_T_1431_data = idxs_T_1431_addr >= 6'h3e ? $random : idxs[idxs_T_1431_addr];
  `endif
  assign idxs_T_1434_addr = {{5'd0}, 1'h1};
  assign idxs_T_1434_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1434_data = idxs[idxs_T_1434_addr];
  `else
  assign idxs_T_1434_data = idxs_T_1434_addr >= 6'h3e ? $random : idxs[idxs_T_1434_addr];
  `endif
  assign idxs_T_1437_addr = {{4'd0}, 2'h2};
  assign idxs_T_1437_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1437_data = idxs[idxs_T_1437_addr];
  `else
  assign idxs_T_1437_data = idxs_T_1437_addr >= 6'h3e ? $random : idxs[idxs_T_1437_addr];
  `endif
  assign idxs_T_1440_addr = {{4'd0}, 2'h3};
  assign idxs_T_1440_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1440_data = idxs[idxs_T_1440_addr];
  `else
  assign idxs_T_1440_data = idxs_T_1440_addr >= 6'h3e ? $random : idxs[idxs_T_1440_addr];
  `endif
  assign idxs_T_1443_addr = {{3'd0}, 3'h4};
  assign idxs_T_1443_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1443_data = idxs[idxs_T_1443_addr];
  `else
  assign idxs_T_1443_data = idxs_T_1443_addr >= 6'h3e ? $random : idxs[idxs_T_1443_addr];
  `endif
  assign idxs_T_1446_addr = {{3'd0}, 3'h5};
  assign idxs_T_1446_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1446_data = idxs[idxs_T_1446_addr];
  `else
  assign idxs_T_1446_data = idxs_T_1446_addr >= 6'h3e ? $random : idxs[idxs_T_1446_addr];
  `endif
  assign idxs_T_1449_addr = {{3'd0}, 3'h6};
  assign idxs_T_1449_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1449_data = idxs[idxs_T_1449_addr];
  `else
  assign idxs_T_1449_data = idxs_T_1449_addr >= 6'h3e ? $random : idxs[idxs_T_1449_addr];
  `endif
  assign idxs_T_1452_addr = {{3'd0}, 3'h7};
  assign idxs_T_1452_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1452_data = idxs[idxs_T_1452_addr];
  `else
  assign idxs_T_1452_data = idxs_T_1452_addr >= 6'h3e ? $random : idxs[idxs_T_1452_addr];
  `endif
  assign idxs_T_1455_addr = {{2'd0}, 4'h8};
  assign idxs_T_1455_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1455_data = idxs[idxs_T_1455_addr];
  `else
  assign idxs_T_1455_data = idxs_T_1455_addr >= 6'h3e ? $random : idxs[idxs_T_1455_addr];
  `endif
  assign idxs_T_1458_addr = {{2'd0}, 4'h9};
  assign idxs_T_1458_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1458_data = idxs[idxs_T_1458_addr];
  `else
  assign idxs_T_1458_data = idxs_T_1458_addr >= 6'h3e ? $random : idxs[idxs_T_1458_addr];
  `endif
  assign idxs_T_1461_addr = {{2'd0}, 4'ha};
  assign idxs_T_1461_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1461_data = idxs[idxs_T_1461_addr];
  `else
  assign idxs_T_1461_data = idxs_T_1461_addr >= 6'h3e ? $random : idxs[idxs_T_1461_addr];
  `endif
  assign idxs_T_1464_addr = {{2'd0}, 4'hb};
  assign idxs_T_1464_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1464_data = idxs[idxs_T_1464_addr];
  `else
  assign idxs_T_1464_data = idxs_T_1464_addr >= 6'h3e ? $random : idxs[idxs_T_1464_addr];
  `endif
  assign idxs_T_1467_addr = {{2'd0}, 4'hc};
  assign idxs_T_1467_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1467_data = idxs[idxs_T_1467_addr];
  `else
  assign idxs_T_1467_data = idxs_T_1467_addr >= 6'h3e ? $random : idxs[idxs_T_1467_addr];
  `endif
  assign idxs_T_1470_addr = {{2'd0}, 4'hd};
  assign idxs_T_1470_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1470_data = idxs[idxs_T_1470_addr];
  `else
  assign idxs_T_1470_data = idxs_T_1470_addr >= 6'h3e ? $random : idxs[idxs_T_1470_addr];
  `endif
  assign idxs_T_1473_addr = {{2'd0}, 4'he};
  assign idxs_T_1473_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1473_data = idxs[idxs_T_1473_addr];
  `else
  assign idxs_T_1473_data = idxs_T_1473_addr >= 6'h3e ? $random : idxs[idxs_T_1473_addr];
  `endif
  assign idxs_T_1476_addr = {{2'd0}, 4'hf};
  assign idxs_T_1476_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1476_data = idxs[idxs_T_1476_addr];
  `else
  assign idxs_T_1476_data = idxs_T_1476_addr >= 6'h3e ? $random : idxs[idxs_T_1476_addr];
  `endif
  assign idxs_T_1479_addr = {{1'd0}, 5'h10};
  assign idxs_T_1479_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1479_data = idxs[idxs_T_1479_addr];
  `else
  assign idxs_T_1479_data = idxs_T_1479_addr >= 6'h3e ? $random : idxs[idxs_T_1479_addr];
  `endif
  assign idxs_T_1482_addr = {{1'd0}, 5'h11};
  assign idxs_T_1482_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1482_data = idxs[idxs_T_1482_addr];
  `else
  assign idxs_T_1482_data = idxs_T_1482_addr >= 6'h3e ? $random : idxs[idxs_T_1482_addr];
  `endif
  assign idxs_T_1485_addr = {{1'd0}, 5'h12};
  assign idxs_T_1485_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1485_data = idxs[idxs_T_1485_addr];
  `else
  assign idxs_T_1485_data = idxs_T_1485_addr >= 6'h3e ? $random : idxs[idxs_T_1485_addr];
  `endif
  assign idxs_T_1488_addr = {{1'd0}, 5'h13};
  assign idxs_T_1488_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1488_data = idxs[idxs_T_1488_addr];
  `else
  assign idxs_T_1488_data = idxs_T_1488_addr >= 6'h3e ? $random : idxs[idxs_T_1488_addr];
  `endif
  assign idxs_T_1491_addr = {{1'd0}, 5'h14};
  assign idxs_T_1491_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1491_data = idxs[idxs_T_1491_addr];
  `else
  assign idxs_T_1491_data = idxs_T_1491_addr >= 6'h3e ? $random : idxs[idxs_T_1491_addr];
  `endif
  assign idxs_T_1494_addr = {{1'd0}, 5'h15};
  assign idxs_T_1494_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1494_data = idxs[idxs_T_1494_addr];
  `else
  assign idxs_T_1494_data = idxs_T_1494_addr >= 6'h3e ? $random : idxs[idxs_T_1494_addr];
  `endif
  assign idxs_T_1497_addr = {{1'd0}, 5'h16};
  assign idxs_T_1497_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1497_data = idxs[idxs_T_1497_addr];
  `else
  assign idxs_T_1497_data = idxs_T_1497_addr >= 6'h3e ? $random : idxs[idxs_T_1497_addr];
  `endif
  assign idxs_T_1500_addr = {{1'd0}, 5'h17};
  assign idxs_T_1500_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1500_data = idxs[idxs_T_1500_addr];
  `else
  assign idxs_T_1500_data = idxs_T_1500_addr >= 6'h3e ? $random : idxs[idxs_T_1500_addr];
  `endif
  assign idxs_T_1503_addr = {{1'd0}, 5'h18};
  assign idxs_T_1503_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1503_data = idxs[idxs_T_1503_addr];
  `else
  assign idxs_T_1503_data = idxs_T_1503_addr >= 6'h3e ? $random : idxs[idxs_T_1503_addr];
  `endif
  assign idxs_T_1506_addr = {{1'd0}, 5'h19};
  assign idxs_T_1506_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1506_data = idxs[idxs_T_1506_addr];
  `else
  assign idxs_T_1506_data = idxs_T_1506_addr >= 6'h3e ? $random : idxs[idxs_T_1506_addr];
  `endif
  assign idxs_T_1509_addr = {{1'd0}, 5'h1a};
  assign idxs_T_1509_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1509_data = idxs[idxs_T_1509_addr];
  `else
  assign idxs_T_1509_data = idxs_T_1509_addr >= 6'h3e ? $random : idxs[idxs_T_1509_addr];
  `endif
  assign idxs_T_1512_addr = {{1'd0}, 5'h1b};
  assign idxs_T_1512_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1512_data = idxs[idxs_T_1512_addr];
  `else
  assign idxs_T_1512_data = idxs_T_1512_addr >= 6'h3e ? $random : idxs[idxs_T_1512_addr];
  `endif
  assign idxs_T_1515_addr = {{1'd0}, 5'h1c};
  assign idxs_T_1515_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1515_data = idxs[idxs_T_1515_addr];
  `else
  assign idxs_T_1515_data = idxs_T_1515_addr >= 6'h3e ? $random : idxs[idxs_T_1515_addr];
  `endif
  assign idxs_T_1518_addr = {{1'd0}, 5'h1d};
  assign idxs_T_1518_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1518_data = idxs[idxs_T_1518_addr];
  `else
  assign idxs_T_1518_data = idxs_T_1518_addr >= 6'h3e ? $random : idxs[idxs_T_1518_addr];
  `endif
  assign idxs_T_1521_addr = {{1'd0}, 5'h1e};
  assign idxs_T_1521_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1521_data = idxs[idxs_T_1521_addr];
  `else
  assign idxs_T_1521_data = idxs_T_1521_addr >= 6'h3e ? $random : idxs[idxs_T_1521_addr];
  `endif
  assign idxs_T_1524_addr = {{1'd0}, 5'h1f};
  assign idxs_T_1524_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1524_data = idxs[idxs_T_1524_addr];
  `else
  assign idxs_T_1524_data = idxs_T_1524_addr >= 6'h3e ? $random : idxs[idxs_T_1524_addr];
  `endif
  assign idxs_T_1527_addr = 6'h20;
  assign idxs_T_1527_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1527_data = idxs[idxs_T_1527_addr];
  `else
  assign idxs_T_1527_data = idxs_T_1527_addr >= 6'h3e ? $random : idxs[idxs_T_1527_addr];
  `endif
  assign idxs_T_1530_addr = 6'h21;
  assign idxs_T_1530_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1530_data = idxs[idxs_T_1530_addr];
  `else
  assign idxs_T_1530_data = idxs_T_1530_addr >= 6'h3e ? $random : idxs[idxs_T_1530_addr];
  `endif
  assign idxs_T_1533_addr = 6'h22;
  assign idxs_T_1533_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1533_data = idxs[idxs_T_1533_addr];
  `else
  assign idxs_T_1533_data = idxs_T_1533_addr >= 6'h3e ? $random : idxs[idxs_T_1533_addr];
  `endif
  assign idxs_T_1536_addr = 6'h23;
  assign idxs_T_1536_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1536_data = idxs[idxs_T_1536_addr];
  `else
  assign idxs_T_1536_data = idxs_T_1536_addr >= 6'h3e ? $random : idxs[idxs_T_1536_addr];
  `endif
  assign idxs_T_1539_addr = 6'h24;
  assign idxs_T_1539_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1539_data = idxs[idxs_T_1539_addr];
  `else
  assign idxs_T_1539_data = idxs_T_1539_addr >= 6'h3e ? $random : idxs[idxs_T_1539_addr];
  `endif
  assign idxs_T_1542_addr = 6'h25;
  assign idxs_T_1542_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1542_data = idxs[idxs_T_1542_addr];
  `else
  assign idxs_T_1542_data = idxs_T_1542_addr >= 6'h3e ? $random : idxs[idxs_T_1542_addr];
  `endif
  assign idxs_T_1545_addr = 6'h26;
  assign idxs_T_1545_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1545_data = idxs[idxs_T_1545_addr];
  `else
  assign idxs_T_1545_data = idxs_T_1545_addr >= 6'h3e ? $random : idxs[idxs_T_1545_addr];
  `endif
  assign idxs_T_1548_addr = 6'h27;
  assign idxs_T_1548_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1548_data = idxs[idxs_T_1548_addr];
  `else
  assign idxs_T_1548_data = idxs_T_1548_addr >= 6'h3e ? $random : idxs[idxs_T_1548_addr];
  `endif
  assign idxs_T_1551_addr = 6'h28;
  assign idxs_T_1551_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1551_data = idxs[idxs_T_1551_addr];
  `else
  assign idxs_T_1551_data = idxs_T_1551_addr >= 6'h3e ? $random : idxs[idxs_T_1551_addr];
  `endif
  assign idxs_T_1554_addr = 6'h29;
  assign idxs_T_1554_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1554_data = idxs[idxs_T_1554_addr];
  `else
  assign idxs_T_1554_data = idxs_T_1554_addr >= 6'h3e ? $random : idxs[idxs_T_1554_addr];
  `endif
  assign idxs_T_1557_addr = 6'h2a;
  assign idxs_T_1557_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1557_data = idxs[idxs_T_1557_addr];
  `else
  assign idxs_T_1557_data = idxs_T_1557_addr >= 6'h3e ? $random : idxs[idxs_T_1557_addr];
  `endif
  assign idxs_T_1560_addr = 6'h2b;
  assign idxs_T_1560_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1560_data = idxs[idxs_T_1560_addr];
  `else
  assign idxs_T_1560_data = idxs_T_1560_addr >= 6'h3e ? $random : idxs[idxs_T_1560_addr];
  `endif
  assign idxs_T_1563_addr = 6'h2c;
  assign idxs_T_1563_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1563_data = idxs[idxs_T_1563_addr];
  `else
  assign idxs_T_1563_data = idxs_T_1563_addr >= 6'h3e ? $random : idxs[idxs_T_1563_addr];
  `endif
  assign idxs_T_1566_addr = 6'h2d;
  assign idxs_T_1566_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1566_data = idxs[idxs_T_1566_addr];
  `else
  assign idxs_T_1566_data = idxs_T_1566_addr >= 6'h3e ? $random : idxs[idxs_T_1566_addr];
  `endif
  assign idxs_T_1569_addr = 6'h2e;
  assign idxs_T_1569_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1569_data = idxs[idxs_T_1569_addr];
  `else
  assign idxs_T_1569_data = idxs_T_1569_addr >= 6'h3e ? $random : idxs[idxs_T_1569_addr];
  `endif
  assign idxs_T_1572_addr = 6'h2f;
  assign idxs_T_1572_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1572_data = idxs[idxs_T_1572_addr];
  `else
  assign idxs_T_1572_data = idxs_T_1572_addr >= 6'h3e ? $random : idxs[idxs_T_1572_addr];
  `endif
  assign idxs_T_1575_addr = 6'h30;
  assign idxs_T_1575_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1575_data = idxs[idxs_T_1575_addr];
  `else
  assign idxs_T_1575_data = idxs_T_1575_addr >= 6'h3e ? $random : idxs[idxs_T_1575_addr];
  `endif
  assign idxs_T_1578_addr = 6'h31;
  assign idxs_T_1578_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1578_data = idxs[idxs_T_1578_addr];
  `else
  assign idxs_T_1578_data = idxs_T_1578_addr >= 6'h3e ? $random : idxs[idxs_T_1578_addr];
  `endif
  assign idxs_T_1581_addr = 6'h32;
  assign idxs_T_1581_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1581_data = idxs[idxs_T_1581_addr];
  `else
  assign idxs_T_1581_data = idxs_T_1581_addr >= 6'h3e ? $random : idxs[idxs_T_1581_addr];
  `endif
  assign idxs_T_1584_addr = 6'h33;
  assign idxs_T_1584_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1584_data = idxs[idxs_T_1584_addr];
  `else
  assign idxs_T_1584_data = idxs_T_1584_addr >= 6'h3e ? $random : idxs[idxs_T_1584_addr];
  `endif
  assign idxs_T_1587_addr = 6'h34;
  assign idxs_T_1587_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1587_data = idxs[idxs_T_1587_addr];
  `else
  assign idxs_T_1587_data = idxs_T_1587_addr >= 6'h3e ? $random : idxs[idxs_T_1587_addr];
  `endif
  assign idxs_T_1590_addr = 6'h35;
  assign idxs_T_1590_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1590_data = idxs[idxs_T_1590_addr];
  `else
  assign idxs_T_1590_data = idxs_T_1590_addr >= 6'h3e ? $random : idxs[idxs_T_1590_addr];
  `endif
  assign idxs_T_1593_addr = 6'h36;
  assign idxs_T_1593_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1593_data = idxs[idxs_T_1593_addr];
  `else
  assign idxs_T_1593_data = idxs_T_1593_addr >= 6'h3e ? $random : idxs[idxs_T_1593_addr];
  `endif
  assign idxs_T_1596_addr = 6'h37;
  assign idxs_T_1596_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1596_data = idxs[idxs_T_1596_addr];
  `else
  assign idxs_T_1596_data = idxs_T_1596_addr >= 6'h3e ? $random : idxs[idxs_T_1596_addr];
  `endif
  assign idxs_T_1599_addr = 6'h38;
  assign idxs_T_1599_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1599_data = idxs[idxs_T_1599_addr];
  `else
  assign idxs_T_1599_data = idxs_T_1599_addr >= 6'h3e ? $random : idxs[idxs_T_1599_addr];
  `endif
  assign idxs_T_1602_addr = 6'h39;
  assign idxs_T_1602_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1602_data = idxs[idxs_T_1602_addr];
  `else
  assign idxs_T_1602_data = idxs_T_1602_addr >= 6'h3e ? $random : idxs[idxs_T_1602_addr];
  `endif
  assign idxs_T_1605_addr = 6'h3a;
  assign idxs_T_1605_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1605_data = idxs[idxs_T_1605_addr];
  `else
  assign idxs_T_1605_data = idxs_T_1605_addr >= 6'h3e ? $random : idxs[idxs_T_1605_addr];
  `endif
  assign idxs_T_1608_addr = 6'h3b;
  assign idxs_T_1608_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1608_data = idxs[idxs_T_1608_addr];
  `else
  assign idxs_T_1608_data = idxs_T_1608_addr >= 6'h3e ? $random : idxs[idxs_T_1608_addr];
  `endif
  assign idxs_T_1611_addr = 6'h3c;
  assign idxs_T_1611_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1611_data = idxs[idxs_T_1611_addr];
  `else
  assign idxs_T_1611_data = idxs_T_1611_addr >= 6'h3e ? $random : idxs[idxs_T_1611_addr];
  `endif
  assign idxs_T_1614_addr = 6'h3d;
  assign idxs_T_1614_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1614_data = idxs[idxs_T_1614_addr];
  `else
  assign idxs_T_1614_data = idxs_T_1614_addr >= 6'h3e ? $random : idxs[idxs_T_1614_addr];
  `endif
  assign idxs_T_1972_addr = {{5'd0}, 1'h0};
  assign idxs_T_1972_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1972_data = idxs[idxs_T_1972_addr];
  `else
  assign idxs_T_1972_data = idxs_T_1972_addr >= 6'h3e ? $random : idxs[idxs_T_1972_addr];
  `endif
  assign idxs_T_1975_addr = {{5'd0}, 1'h1};
  assign idxs_T_1975_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1975_data = idxs[idxs_T_1975_addr];
  `else
  assign idxs_T_1975_data = idxs_T_1975_addr >= 6'h3e ? $random : idxs[idxs_T_1975_addr];
  `endif
  assign idxs_T_1978_addr = {{4'd0}, 2'h2};
  assign idxs_T_1978_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1978_data = idxs[idxs_T_1978_addr];
  `else
  assign idxs_T_1978_data = idxs_T_1978_addr >= 6'h3e ? $random : idxs[idxs_T_1978_addr];
  `endif
  assign idxs_T_1981_addr = {{4'd0}, 2'h3};
  assign idxs_T_1981_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1981_data = idxs[idxs_T_1981_addr];
  `else
  assign idxs_T_1981_data = idxs_T_1981_addr >= 6'h3e ? $random : idxs[idxs_T_1981_addr];
  `endif
  assign idxs_T_1984_addr = {{3'd0}, 3'h4};
  assign idxs_T_1984_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1984_data = idxs[idxs_T_1984_addr];
  `else
  assign idxs_T_1984_data = idxs_T_1984_addr >= 6'h3e ? $random : idxs[idxs_T_1984_addr];
  `endif
  assign idxs_T_1987_addr = {{3'd0}, 3'h5};
  assign idxs_T_1987_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1987_data = idxs[idxs_T_1987_addr];
  `else
  assign idxs_T_1987_data = idxs_T_1987_addr >= 6'h3e ? $random : idxs[idxs_T_1987_addr];
  `endif
  assign idxs_T_1990_addr = {{3'd0}, 3'h6};
  assign idxs_T_1990_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1990_data = idxs[idxs_T_1990_addr];
  `else
  assign idxs_T_1990_data = idxs_T_1990_addr >= 6'h3e ? $random : idxs[idxs_T_1990_addr];
  `endif
  assign idxs_T_1993_addr = {{3'd0}, 3'h7};
  assign idxs_T_1993_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1993_data = idxs[idxs_T_1993_addr];
  `else
  assign idxs_T_1993_data = idxs_T_1993_addr >= 6'h3e ? $random : idxs[idxs_T_1993_addr];
  `endif
  assign idxs_T_1996_addr = {{2'd0}, 4'h8};
  assign idxs_T_1996_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1996_data = idxs[idxs_T_1996_addr];
  `else
  assign idxs_T_1996_data = idxs_T_1996_addr >= 6'h3e ? $random : idxs[idxs_T_1996_addr];
  `endif
  assign idxs_T_1999_addr = {{2'd0}, 4'h9};
  assign idxs_T_1999_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1999_data = idxs[idxs_T_1999_addr];
  `else
  assign idxs_T_1999_data = idxs_T_1999_addr >= 6'h3e ? $random : idxs[idxs_T_1999_addr];
  `endif
  assign idxs_T_2002_addr = {{2'd0}, 4'ha};
  assign idxs_T_2002_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2002_data = idxs[idxs_T_2002_addr];
  `else
  assign idxs_T_2002_data = idxs_T_2002_addr >= 6'h3e ? $random : idxs[idxs_T_2002_addr];
  `endif
  assign idxs_T_2005_addr = {{2'd0}, 4'hb};
  assign idxs_T_2005_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2005_data = idxs[idxs_T_2005_addr];
  `else
  assign idxs_T_2005_data = idxs_T_2005_addr >= 6'h3e ? $random : idxs[idxs_T_2005_addr];
  `endif
  assign idxs_T_2008_addr = {{2'd0}, 4'hc};
  assign idxs_T_2008_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2008_data = idxs[idxs_T_2008_addr];
  `else
  assign idxs_T_2008_data = idxs_T_2008_addr >= 6'h3e ? $random : idxs[idxs_T_2008_addr];
  `endif
  assign idxs_T_2011_addr = {{2'd0}, 4'hd};
  assign idxs_T_2011_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2011_data = idxs[idxs_T_2011_addr];
  `else
  assign idxs_T_2011_data = idxs_T_2011_addr >= 6'h3e ? $random : idxs[idxs_T_2011_addr];
  `endif
  assign idxs_T_2014_addr = {{2'd0}, 4'he};
  assign idxs_T_2014_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2014_data = idxs[idxs_T_2014_addr];
  `else
  assign idxs_T_2014_data = idxs_T_2014_addr >= 6'h3e ? $random : idxs[idxs_T_2014_addr];
  `endif
  assign idxs_T_2017_addr = {{2'd0}, 4'hf};
  assign idxs_T_2017_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2017_data = idxs[idxs_T_2017_addr];
  `else
  assign idxs_T_2017_data = idxs_T_2017_addr >= 6'h3e ? $random : idxs[idxs_T_2017_addr];
  `endif
  assign idxs_T_2020_addr = {{1'd0}, 5'h10};
  assign idxs_T_2020_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2020_data = idxs[idxs_T_2020_addr];
  `else
  assign idxs_T_2020_data = idxs_T_2020_addr >= 6'h3e ? $random : idxs[idxs_T_2020_addr];
  `endif
  assign idxs_T_2023_addr = {{1'd0}, 5'h11};
  assign idxs_T_2023_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2023_data = idxs[idxs_T_2023_addr];
  `else
  assign idxs_T_2023_data = idxs_T_2023_addr >= 6'h3e ? $random : idxs[idxs_T_2023_addr];
  `endif
  assign idxs_T_2026_addr = {{1'd0}, 5'h12};
  assign idxs_T_2026_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2026_data = idxs[idxs_T_2026_addr];
  `else
  assign idxs_T_2026_data = idxs_T_2026_addr >= 6'h3e ? $random : idxs[idxs_T_2026_addr];
  `endif
  assign idxs_T_2029_addr = {{1'd0}, 5'h13};
  assign idxs_T_2029_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2029_data = idxs[idxs_T_2029_addr];
  `else
  assign idxs_T_2029_data = idxs_T_2029_addr >= 6'h3e ? $random : idxs[idxs_T_2029_addr];
  `endif
  assign idxs_T_2032_addr = {{1'd0}, 5'h14};
  assign idxs_T_2032_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2032_data = idxs[idxs_T_2032_addr];
  `else
  assign idxs_T_2032_data = idxs_T_2032_addr >= 6'h3e ? $random : idxs[idxs_T_2032_addr];
  `endif
  assign idxs_T_2035_addr = {{1'd0}, 5'h15};
  assign idxs_T_2035_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2035_data = idxs[idxs_T_2035_addr];
  `else
  assign idxs_T_2035_data = idxs_T_2035_addr >= 6'h3e ? $random : idxs[idxs_T_2035_addr];
  `endif
  assign idxs_T_2038_addr = {{1'd0}, 5'h16};
  assign idxs_T_2038_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2038_data = idxs[idxs_T_2038_addr];
  `else
  assign idxs_T_2038_data = idxs_T_2038_addr >= 6'h3e ? $random : idxs[idxs_T_2038_addr];
  `endif
  assign idxs_T_2041_addr = {{1'd0}, 5'h17};
  assign idxs_T_2041_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2041_data = idxs[idxs_T_2041_addr];
  `else
  assign idxs_T_2041_data = idxs_T_2041_addr >= 6'h3e ? $random : idxs[idxs_T_2041_addr];
  `endif
  assign idxs_T_2044_addr = {{1'd0}, 5'h18};
  assign idxs_T_2044_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2044_data = idxs[idxs_T_2044_addr];
  `else
  assign idxs_T_2044_data = idxs_T_2044_addr >= 6'h3e ? $random : idxs[idxs_T_2044_addr];
  `endif
  assign idxs_T_2047_addr = {{1'd0}, 5'h19};
  assign idxs_T_2047_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2047_data = idxs[idxs_T_2047_addr];
  `else
  assign idxs_T_2047_data = idxs_T_2047_addr >= 6'h3e ? $random : idxs[idxs_T_2047_addr];
  `endif
  assign idxs_T_2050_addr = {{1'd0}, 5'h1a};
  assign idxs_T_2050_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2050_data = idxs[idxs_T_2050_addr];
  `else
  assign idxs_T_2050_data = idxs_T_2050_addr >= 6'h3e ? $random : idxs[idxs_T_2050_addr];
  `endif
  assign idxs_T_2053_addr = {{1'd0}, 5'h1b};
  assign idxs_T_2053_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2053_data = idxs[idxs_T_2053_addr];
  `else
  assign idxs_T_2053_data = idxs_T_2053_addr >= 6'h3e ? $random : idxs[idxs_T_2053_addr];
  `endif
  assign idxs_T_2056_addr = {{1'd0}, 5'h1c};
  assign idxs_T_2056_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2056_data = idxs[idxs_T_2056_addr];
  `else
  assign idxs_T_2056_data = idxs_T_2056_addr >= 6'h3e ? $random : idxs[idxs_T_2056_addr];
  `endif
  assign idxs_T_2059_addr = {{1'd0}, 5'h1d};
  assign idxs_T_2059_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2059_data = idxs[idxs_T_2059_addr];
  `else
  assign idxs_T_2059_data = idxs_T_2059_addr >= 6'h3e ? $random : idxs[idxs_T_2059_addr];
  `endif
  assign idxs_T_2062_addr = {{1'd0}, 5'h1e};
  assign idxs_T_2062_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2062_data = idxs[idxs_T_2062_addr];
  `else
  assign idxs_T_2062_data = idxs_T_2062_addr >= 6'h3e ? $random : idxs[idxs_T_2062_addr];
  `endif
  assign idxs_T_2065_addr = {{1'd0}, 5'h1f};
  assign idxs_T_2065_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2065_data = idxs[idxs_T_2065_addr];
  `else
  assign idxs_T_2065_data = idxs_T_2065_addr >= 6'h3e ? $random : idxs[idxs_T_2065_addr];
  `endif
  assign idxs_T_2068_addr = 6'h20;
  assign idxs_T_2068_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2068_data = idxs[idxs_T_2068_addr];
  `else
  assign idxs_T_2068_data = idxs_T_2068_addr >= 6'h3e ? $random : idxs[idxs_T_2068_addr];
  `endif
  assign idxs_T_2071_addr = 6'h21;
  assign idxs_T_2071_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2071_data = idxs[idxs_T_2071_addr];
  `else
  assign idxs_T_2071_data = idxs_T_2071_addr >= 6'h3e ? $random : idxs[idxs_T_2071_addr];
  `endif
  assign idxs_T_2074_addr = 6'h22;
  assign idxs_T_2074_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2074_data = idxs[idxs_T_2074_addr];
  `else
  assign idxs_T_2074_data = idxs_T_2074_addr >= 6'h3e ? $random : idxs[idxs_T_2074_addr];
  `endif
  assign idxs_T_2077_addr = 6'h23;
  assign idxs_T_2077_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2077_data = idxs[idxs_T_2077_addr];
  `else
  assign idxs_T_2077_data = idxs_T_2077_addr >= 6'h3e ? $random : idxs[idxs_T_2077_addr];
  `endif
  assign idxs_T_2080_addr = 6'h24;
  assign idxs_T_2080_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2080_data = idxs[idxs_T_2080_addr];
  `else
  assign idxs_T_2080_data = idxs_T_2080_addr >= 6'h3e ? $random : idxs[idxs_T_2080_addr];
  `endif
  assign idxs_T_2083_addr = 6'h25;
  assign idxs_T_2083_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2083_data = idxs[idxs_T_2083_addr];
  `else
  assign idxs_T_2083_data = idxs_T_2083_addr >= 6'h3e ? $random : idxs[idxs_T_2083_addr];
  `endif
  assign idxs_T_2086_addr = 6'h26;
  assign idxs_T_2086_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2086_data = idxs[idxs_T_2086_addr];
  `else
  assign idxs_T_2086_data = idxs_T_2086_addr >= 6'h3e ? $random : idxs[idxs_T_2086_addr];
  `endif
  assign idxs_T_2089_addr = 6'h27;
  assign idxs_T_2089_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2089_data = idxs[idxs_T_2089_addr];
  `else
  assign idxs_T_2089_data = idxs_T_2089_addr >= 6'h3e ? $random : idxs[idxs_T_2089_addr];
  `endif
  assign idxs_T_2092_addr = 6'h28;
  assign idxs_T_2092_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2092_data = idxs[idxs_T_2092_addr];
  `else
  assign idxs_T_2092_data = idxs_T_2092_addr >= 6'h3e ? $random : idxs[idxs_T_2092_addr];
  `endif
  assign idxs_T_2095_addr = 6'h29;
  assign idxs_T_2095_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2095_data = idxs[idxs_T_2095_addr];
  `else
  assign idxs_T_2095_data = idxs_T_2095_addr >= 6'h3e ? $random : idxs[idxs_T_2095_addr];
  `endif
  assign idxs_T_2098_addr = 6'h2a;
  assign idxs_T_2098_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2098_data = idxs[idxs_T_2098_addr];
  `else
  assign idxs_T_2098_data = idxs_T_2098_addr >= 6'h3e ? $random : idxs[idxs_T_2098_addr];
  `endif
  assign idxs_T_2101_addr = 6'h2b;
  assign idxs_T_2101_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2101_data = idxs[idxs_T_2101_addr];
  `else
  assign idxs_T_2101_data = idxs_T_2101_addr >= 6'h3e ? $random : idxs[idxs_T_2101_addr];
  `endif
  assign idxs_T_2104_addr = 6'h2c;
  assign idxs_T_2104_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2104_data = idxs[idxs_T_2104_addr];
  `else
  assign idxs_T_2104_data = idxs_T_2104_addr >= 6'h3e ? $random : idxs[idxs_T_2104_addr];
  `endif
  assign idxs_T_2107_addr = 6'h2d;
  assign idxs_T_2107_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2107_data = idxs[idxs_T_2107_addr];
  `else
  assign idxs_T_2107_data = idxs_T_2107_addr >= 6'h3e ? $random : idxs[idxs_T_2107_addr];
  `endif
  assign idxs_T_2110_addr = 6'h2e;
  assign idxs_T_2110_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2110_data = idxs[idxs_T_2110_addr];
  `else
  assign idxs_T_2110_data = idxs_T_2110_addr >= 6'h3e ? $random : idxs[idxs_T_2110_addr];
  `endif
  assign idxs_T_2113_addr = 6'h2f;
  assign idxs_T_2113_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2113_data = idxs[idxs_T_2113_addr];
  `else
  assign idxs_T_2113_data = idxs_T_2113_addr >= 6'h3e ? $random : idxs[idxs_T_2113_addr];
  `endif
  assign idxs_T_2116_addr = 6'h30;
  assign idxs_T_2116_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2116_data = idxs[idxs_T_2116_addr];
  `else
  assign idxs_T_2116_data = idxs_T_2116_addr >= 6'h3e ? $random : idxs[idxs_T_2116_addr];
  `endif
  assign idxs_T_2119_addr = 6'h31;
  assign idxs_T_2119_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2119_data = idxs[idxs_T_2119_addr];
  `else
  assign idxs_T_2119_data = idxs_T_2119_addr >= 6'h3e ? $random : idxs[idxs_T_2119_addr];
  `endif
  assign idxs_T_2122_addr = 6'h32;
  assign idxs_T_2122_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2122_data = idxs[idxs_T_2122_addr];
  `else
  assign idxs_T_2122_data = idxs_T_2122_addr >= 6'h3e ? $random : idxs[idxs_T_2122_addr];
  `endif
  assign idxs_T_2125_addr = 6'h33;
  assign idxs_T_2125_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2125_data = idxs[idxs_T_2125_addr];
  `else
  assign idxs_T_2125_data = idxs_T_2125_addr >= 6'h3e ? $random : idxs[idxs_T_2125_addr];
  `endif
  assign idxs_T_2128_addr = 6'h34;
  assign idxs_T_2128_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2128_data = idxs[idxs_T_2128_addr];
  `else
  assign idxs_T_2128_data = idxs_T_2128_addr >= 6'h3e ? $random : idxs[idxs_T_2128_addr];
  `endif
  assign idxs_T_2131_addr = 6'h35;
  assign idxs_T_2131_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2131_data = idxs[idxs_T_2131_addr];
  `else
  assign idxs_T_2131_data = idxs_T_2131_addr >= 6'h3e ? $random : idxs[idxs_T_2131_addr];
  `endif
  assign idxs_T_2134_addr = 6'h36;
  assign idxs_T_2134_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2134_data = idxs[idxs_T_2134_addr];
  `else
  assign idxs_T_2134_data = idxs_T_2134_addr >= 6'h3e ? $random : idxs[idxs_T_2134_addr];
  `endif
  assign idxs_T_2137_addr = 6'h37;
  assign idxs_T_2137_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2137_data = idxs[idxs_T_2137_addr];
  `else
  assign idxs_T_2137_data = idxs_T_2137_addr >= 6'h3e ? $random : idxs[idxs_T_2137_addr];
  `endif
  assign idxs_T_2140_addr = 6'h38;
  assign idxs_T_2140_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2140_data = idxs[idxs_T_2140_addr];
  `else
  assign idxs_T_2140_data = idxs_T_2140_addr >= 6'h3e ? $random : idxs[idxs_T_2140_addr];
  `endif
  assign idxs_T_2143_addr = 6'h39;
  assign idxs_T_2143_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2143_data = idxs[idxs_T_2143_addr];
  `else
  assign idxs_T_2143_data = idxs_T_2143_addr >= 6'h3e ? $random : idxs[idxs_T_2143_addr];
  `endif
  assign idxs_T_2146_addr = 6'h3a;
  assign idxs_T_2146_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2146_data = idxs[idxs_T_2146_addr];
  `else
  assign idxs_T_2146_data = idxs_T_2146_addr >= 6'h3e ? $random : idxs[idxs_T_2146_addr];
  `endif
  assign idxs_T_2149_addr = 6'h3b;
  assign idxs_T_2149_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2149_data = idxs[idxs_T_2149_addr];
  `else
  assign idxs_T_2149_data = idxs_T_2149_addr >= 6'h3e ? $random : idxs[idxs_T_2149_addr];
  `endif
  assign idxs_T_2152_addr = 6'h3c;
  assign idxs_T_2152_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2152_data = idxs[idxs_T_2152_addr];
  `else
  assign idxs_T_2152_data = idxs_T_2152_addr >= 6'h3e ? $random : idxs[idxs_T_2152_addr];
  `endif
  assign idxs_T_2155_addr = 6'h3d;
  assign idxs_T_2155_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2155_data = idxs[idxs_T_2155_addr];
  `else
  assign idxs_T_2155_data = idxs_T_2155_addr >= 6'h3e ? $random : idxs[idxs_T_2155_addr];
  `endif
  assign idxs_T_2872_data = r_btb_update_bits_pc[11:0];
  assign idxs_T_2872_addr = T_2550;
  assign idxs_T_2872_mask = r_btb_update_valid;
  assign idxs_T_2872_en = r_btb_update_valid;
  assign idxPages_T_578_addr = {{5'd0}, 1'h0};
  assign idxPages_T_578_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_578_data = idxPages[idxPages_T_578_addr];
  `else
  assign idxPages_T_578_data = idxPages_T_578_addr >= 6'h3e ? $random : idxPages[idxPages_T_578_addr];
  `endif
  assign idxPages_T_583_addr = {{5'd0}, 1'h1};
  assign idxPages_T_583_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_583_data = idxPages[idxPages_T_583_addr];
  `else
  assign idxPages_T_583_data = idxPages_T_583_addr >= 6'h3e ? $random : idxPages[idxPages_T_583_addr];
  `endif
  assign idxPages_T_588_addr = {{4'd0}, 2'h2};
  assign idxPages_T_588_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_588_data = idxPages[idxPages_T_588_addr];
  `else
  assign idxPages_T_588_data = idxPages_T_588_addr >= 6'h3e ? $random : idxPages[idxPages_T_588_addr];
  `endif
  assign idxPages_T_593_addr = {{4'd0}, 2'h3};
  assign idxPages_T_593_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_593_data = idxPages[idxPages_T_593_addr];
  `else
  assign idxPages_T_593_data = idxPages_T_593_addr >= 6'h3e ? $random : idxPages[idxPages_T_593_addr];
  `endif
  assign idxPages_T_598_addr = {{3'd0}, 3'h4};
  assign idxPages_T_598_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_598_data = idxPages[idxPages_T_598_addr];
  `else
  assign idxPages_T_598_data = idxPages_T_598_addr >= 6'h3e ? $random : idxPages[idxPages_T_598_addr];
  `endif
  assign idxPages_T_603_addr = {{3'd0}, 3'h5};
  assign idxPages_T_603_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_603_data = idxPages[idxPages_T_603_addr];
  `else
  assign idxPages_T_603_data = idxPages_T_603_addr >= 6'h3e ? $random : idxPages[idxPages_T_603_addr];
  `endif
  assign idxPages_T_608_addr = {{3'd0}, 3'h6};
  assign idxPages_T_608_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_608_data = idxPages[idxPages_T_608_addr];
  `else
  assign idxPages_T_608_data = idxPages_T_608_addr >= 6'h3e ? $random : idxPages[idxPages_T_608_addr];
  `endif
  assign idxPages_T_613_addr = {{3'd0}, 3'h7};
  assign idxPages_T_613_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_613_data = idxPages[idxPages_T_613_addr];
  `else
  assign idxPages_T_613_data = idxPages_T_613_addr >= 6'h3e ? $random : idxPages[idxPages_T_613_addr];
  `endif
  assign idxPages_T_618_addr = {{2'd0}, 4'h8};
  assign idxPages_T_618_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_618_data = idxPages[idxPages_T_618_addr];
  `else
  assign idxPages_T_618_data = idxPages_T_618_addr >= 6'h3e ? $random : idxPages[idxPages_T_618_addr];
  `endif
  assign idxPages_T_623_addr = {{2'd0}, 4'h9};
  assign idxPages_T_623_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_623_data = idxPages[idxPages_T_623_addr];
  `else
  assign idxPages_T_623_data = idxPages_T_623_addr >= 6'h3e ? $random : idxPages[idxPages_T_623_addr];
  `endif
  assign idxPages_T_628_addr = {{2'd0}, 4'ha};
  assign idxPages_T_628_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_628_data = idxPages[idxPages_T_628_addr];
  `else
  assign idxPages_T_628_data = idxPages_T_628_addr >= 6'h3e ? $random : idxPages[idxPages_T_628_addr];
  `endif
  assign idxPages_T_633_addr = {{2'd0}, 4'hb};
  assign idxPages_T_633_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_633_data = idxPages[idxPages_T_633_addr];
  `else
  assign idxPages_T_633_data = idxPages_T_633_addr >= 6'h3e ? $random : idxPages[idxPages_T_633_addr];
  `endif
  assign idxPages_T_638_addr = {{2'd0}, 4'hc};
  assign idxPages_T_638_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_638_data = idxPages[idxPages_T_638_addr];
  `else
  assign idxPages_T_638_data = idxPages_T_638_addr >= 6'h3e ? $random : idxPages[idxPages_T_638_addr];
  `endif
  assign idxPages_T_643_addr = {{2'd0}, 4'hd};
  assign idxPages_T_643_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_643_data = idxPages[idxPages_T_643_addr];
  `else
  assign idxPages_T_643_data = idxPages_T_643_addr >= 6'h3e ? $random : idxPages[idxPages_T_643_addr];
  `endif
  assign idxPages_T_648_addr = {{2'd0}, 4'he};
  assign idxPages_T_648_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_648_data = idxPages[idxPages_T_648_addr];
  `else
  assign idxPages_T_648_data = idxPages_T_648_addr >= 6'h3e ? $random : idxPages[idxPages_T_648_addr];
  `endif
  assign idxPages_T_653_addr = {{2'd0}, 4'hf};
  assign idxPages_T_653_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_653_data = idxPages[idxPages_T_653_addr];
  `else
  assign idxPages_T_653_data = idxPages_T_653_addr >= 6'h3e ? $random : idxPages[idxPages_T_653_addr];
  `endif
  assign idxPages_T_658_addr = {{1'd0}, 5'h10};
  assign idxPages_T_658_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_658_data = idxPages[idxPages_T_658_addr];
  `else
  assign idxPages_T_658_data = idxPages_T_658_addr >= 6'h3e ? $random : idxPages[idxPages_T_658_addr];
  `endif
  assign idxPages_T_663_addr = {{1'd0}, 5'h11};
  assign idxPages_T_663_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_663_data = idxPages[idxPages_T_663_addr];
  `else
  assign idxPages_T_663_data = idxPages_T_663_addr >= 6'h3e ? $random : idxPages[idxPages_T_663_addr];
  `endif
  assign idxPages_T_668_addr = {{1'd0}, 5'h12};
  assign idxPages_T_668_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_668_data = idxPages[idxPages_T_668_addr];
  `else
  assign idxPages_T_668_data = idxPages_T_668_addr >= 6'h3e ? $random : idxPages[idxPages_T_668_addr];
  `endif
  assign idxPages_T_673_addr = {{1'd0}, 5'h13};
  assign idxPages_T_673_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_673_data = idxPages[idxPages_T_673_addr];
  `else
  assign idxPages_T_673_data = idxPages_T_673_addr >= 6'h3e ? $random : idxPages[idxPages_T_673_addr];
  `endif
  assign idxPages_T_678_addr = {{1'd0}, 5'h14};
  assign idxPages_T_678_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_678_data = idxPages[idxPages_T_678_addr];
  `else
  assign idxPages_T_678_data = idxPages_T_678_addr >= 6'h3e ? $random : idxPages[idxPages_T_678_addr];
  `endif
  assign idxPages_T_683_addr = {{1'd0}, 5'h15};
  assign idxPages_T_683_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_683_data = idxPages[idxPages_T_683_addr];
  `else
  assign idxPages_T_683_data = idxPages_T_683_addr >= 6'h3e ? $random : idxPages[idxPages_T_683_addr];
  `endif
  assign idxPages_T_688_addr = {{1'd0}, 5'h16};
  assign idxPages_T_688_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_688_data = idxPages[idxPages_T_688_addr];
  `else
  assign idxPages_T_688_data = idxPages_T_688_addr >= 6'h3e ? $random : idxPages[idxPages_T_688_addr];
  `endif
  assign idxPages_T_693_addr = {{1'd0}, 5'h17};
  assign idxPages_T_693_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_693_data = idxPages[idxPages_T_693_addr];
  `else
  assign idxPages_T_693_data = idxPages_T_693_addr >= 6'h3e ? $random : idxPages[idxPages_T_693_addr];
  `endif
  assign idxPages_T_698_addr = {{1'd0}, 5'h18};
  assign idxPages_T_698_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_698_data = idxPages[idxPages_T_698_addr];
  `else
  assign idxPages_T_698_data = idxPages_T_698_addr >= 6'h3e ? $random : idxPages[idxPages_T_698_addr];
  `endif
  assign idxPages_T_703_addr = {{1'd0}, 5'h19};
  assign idxPages_T_703_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_703_data = idxPages[idxPages_T_703_addr];
  `else
  assign idxPages_T_703_data = idxPages_T_703_addr >= 6'h3e ? $random : idxPages[idxPages_T_703_addr];
  `endif
  assign idxPages_T_708_addr = {{1'd0}, 5'h1a};
  assign idxPages_T_708_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_708_data = idxPages[idxPages_T_708_addr];
  `else
  assign idxPages_T_708_data = idxPages_T_708_addr >= 6'h3e ? $random : idxPages[idxPages_T_708_addr];
  `endif
  assign idxPages_T_713_addr = {{1'd0}, 5'h1b};
  assign idxPages_T_713_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_713_data = idxPages[idxPages_T_713_addr];
  `else
  assign idxPages_T_713_data = idxPages_T_713_addr >= 6'h3e ? $random : idxPages[idxPages_T_713_addr];
  `endif
  assign idxPages_T_718_addr = {{1'd0}, 5'h1c};
  assign idxPages_T_718_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_718_data = idxPages[idxPages_T_718_addr];
  `else
  assign idxPages_T_718_data = idxPages_T_718_addr >= 6'h3e ? $random : idxPages[idxPages_T_718_addr];
  `endif
  assign idxPages_T_723_addr = {{1'd0}, 5'h1d};
  assign idxPages_T_723_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_723_data = idxPages[idxPages_T_723_addr];
  `else
  assign idxPages_T_723_data = idxPages_T_723_addr >= 6'h3e ? $random : idxPages[idxPages_T_723_addr];
  `endif
  assign idxPages_T_728_addr = {{1'd0}, 5'h1e};
  assign idxPages_T_728_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_728_data = idxPages[idxPages_T_728_addr];
  `else
  assign idxPages_T_728_data = idxPages_T_728_addr >= 6'h3e ? $random : idxPages[idxPages_T_728_addr];
  `endif
  assign idxPages_T_733_addr = {{1'd0}, 5'h1f};
  assign idxPages_T_733_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_733_data = idxPages[idxPages_T_733_addr];
  `else
  assign idxPages_T_733_data = idxPages_T_733_addr >= 6'h3e ? $random : idxPages[idxPages_T_733_addr];
  `endif
  assign idxPages_T_738_addr = 6'h20;
  assign idxPages_T_738_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_738_data = idxPages[idxPages_T_738_addr];
  `else
  assign idxPages_T_738_data = idxPages_T_738_addr >= 6'h3e ? $random : idxPages[idxPages_T_738_addr];
  `endif
  assign idxPages_T_743_addr = 6'h21;
  assign idxPages_T_743_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_743_data = idxPages[idxPages_T_743_addr];
  `else
  assign idxPages_T_743_data = idxPages_T_743_addr >= 6'h3e ? $random : idxPages[idxPages_T_743_addr];
  `endif
  assign idxPages_T_748_addr = 6'h22;
  assign idxPages_T_748_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_748_data = idxPages[idxPages_T_748_addr];
  `else
  assign idxPages_T_748_data = idxPages_T_748_addr >= 6'h3e ? $random : idxPages[idxPages_T_748_addr];
  `endif
  assign idxPages_T_753_addr = 6'h23;
  assign idxPages_T_753_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_753_data = idxPages[idxPages_T_753_addr];
  `else
  assign idxPages_T_753_data = idxPages_T_753_addr >= 6'h3e ? $random : idxPages[idxPages_T_753_addr];
  `endif
  assign idxPages_T_758_addr = 6'h24;
  assign idxPages_T_758_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_758_data = idxPages[idxPages_T_758_addr];
  `else
  assign idxPages_T_758_data = idxPages_T_758_addr >= 6'h3e ? $random : idxPages[idxPages_T_758_addr];
  `endif
  assign idxPages_T_763_addr = 6'h25;
  assign idxPages_T_763_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_763_data = idxPages[idxPages_T_763_addr];
  `else
  assign idxPages_T_763_data = idxPages_T_763_addr >= 6'h3e ? $random : idxPages[idxPages_T_763_addr];
  `endif
  assign idxPages_T_768_addr = 6'h26;
  assign idxPages_T_768_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_768_data = idxPages[idxPages_T_768_addr];
  `else
  assign idxPages_T_768_data = idxPages_T_768_addr >= 6'h3e ? $random : idxPages[idxPages_T_768_addr];
  `endif
  assign idxPages_T_773_addr = 6'h27;
  assign idxPages_T_773_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_773_data = idxPages[idxPages_T_773_addr];
  `else
  assign idxPages_T_773_data = idxPages_T_773_addr >= 6'h3e ? $random : idxPages[idxPages_T_773_addr];
  `endif
  assign idxPages_T_778_addr = 6'h28;
  assign idxPages_T_778_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_778_data = idxPages[idxPages_T_778_addr];
  `else
  assign idxPages_T_778_data = idxPages_T_778_addr >= 6'h3e ? $random : idxPages[idxPages_T_778_addr];
  `endif
  assign idxPages_T_783_addr = 6'h29;
  assign idxPages_T_783_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_783_data = idxPages[idxPages_T_783_addr];
  `else
  assign idxPages_T_783_data = idxPages_T_783_addr >= 6'h3e ? $random : idxPages[idxPages_T_783_addr];
  `endif
  assign idxPages_T_788_addr = 6'h2a;
  assign idxPages_T_788_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_788_data = idxPages[idxPages_T_788_addr];
  `else
  assign idxPages_T_788_data = idxPages_T_788_addr >= 6'h3e ? $random : idxPages[idxPages_T_788_addr];
  `endif
  assign idxPages_T_793_addr = 6'h2b;
  assign idxPages_T_793_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_793_data = idxPages[idxPages_T_793_addr];
  `else
  assign idxPages_T_793_data = idxPages_T_793_addr >= 6'h3e ? $random : idxPages[idxPages_T_793_addr];
  `endif
  assign idxPages_T_798_addr = 6'h2c;
  assign idxPages_T_798_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_798_data = idxPages[idxPages_T_798_addr];
  `else
  assign idxPages_T_798_data = idxPages_T_798_addr >= 6'h3e ? $random : idxPages[idxPages_T_798_addr];
  `endif
  assign idxPages_T_803_addr = 6'h2d;
  assign idxPages_T_803_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_803_data = idxPages[idxPages_T_803_addr];
  `else
  assign idxPages_T_803_data = idxPages_T_803_addr >= 6'h3e ? $random : idxPages[idxPages_T_803_addr];
  `endif
  assign idxPages_T_808_addr = 6'h2e;
  assign idxPages_T_808_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_808_data = idxPages[idxPages_T_808_addr];
  `else
  assign idxPages_T_808_data = idxPages_T_808_addr >= 6'h3e ? $random : idxPages[idxPages_T_808_addr];
  `endif
  assign idxPages_T_813_addr = 6'h2f;
  assign idxPages_T_813_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_813_data = idxPages[idxPages_T_813_addr];
  `else
  assign idxPages_T_813_data = idxPages_T_813_addr >= 6'h3e ? $random : idxPages[idxPages_T_813_addr];
  `endif
  assign idxPages_T_818_addr = 6'h30;
  assign idxPages_T_818_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_818_data = idxPages[idxPages_T_818_addr];
  `else
  assign idxPages_T_818_data = idxPages_T_818_addr >= 6'h3e ? $random : idxPages[idxPages_T_818_addr];
  `endif
  assign idxPages_T_823_addr = 6'h31;
  assign idxPages_T_823_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_823_data = idxPages[idxPages_T_823_addr];
  `else
  assign idxPages_T_823_data = idxPages_T_823_addr >= 6'h3e ? $random : idxPages[idxPages_T_823_addr];
  `endif
  assign idxPages_T_828_addr = 6'h32;
  assign idxPages_T_828_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_828_data = idxPages[idxPages_T_828_addr];
  `else
  assign idxPages_T_828_data = idxPages_T_828_addr >= 6'h3e ? $random : idxPages[idxPages_T_828_addr];
  `endif
  assign idxPages_T_833_addr = 6'h33;
  assign idxPages_T_833_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_833_data = idxPages[idxPages_T_833_addr];
  `else
  assign idxPages_T_833_data = idxPages_T_833_addr >= 6'h3e ? $random : idxPages[idxPages_T_833_addr];
  `endif
  assign idxPages_T_838_addr = 6'h34;
  assign idxPages_T_838_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_838_data = idxPages[idxPages_T_838_addr];
  `else
  assign idxPages_T_838_data = idxPages_T_838_addr >= 6'h3e ? $random : idxPages[idxPages_T_838_addr];
  `endif
  assign idxPages_T_843_addr = 6'h35;
  assign idxPages_T_843_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_843_data = idxPages[idxPages_T_843_addr];
  `else
  assign idxPages_T_843_data = idxPages_T_843_addr >= 6'h3e ? $random : idxPages[idxPages_T_843_addr];
  `endif
  assign idxPages_T_848_addr = 6'h36;
  assign idxPages_T_848_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_848_data = idxPages[idxPages_T_848_addr];
  `else
  assign idxPages_T_848_data = idxPages_T_848_addr >= 6'h3e ? $random : idxPages[idxPages_T_848_addr];
  `endif
  assign idxPages_T_853_addr = 6'h37;
  assign idxPages_T_853_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_853_data = idxPages[idxPages_T_853_addr];
  `else
  assign idxPages_T_853_data = idxPages_T_853_addr >= 6'h3e ? $random : idxPages[idxPages_T_853_addr];
  `endif
  assign idxPages_T_858_addr = 6'h38;
  assign idxPages_T_858_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_858_data = idxPages[idxPages_T_858_addr];
  `else
  assign idxPages_T_858_data = idxPages_T_858_addr >= 6'h3e ? $random : idxPages[idxPages_T_858_addr];
  `endif
  assign idxPages_T_863_addr = 6'h39;
  assign idxPages_T_863_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_863_data = idxPages[idxPages_T_863_addr];
  `else
  assign idxPages_T_863_data = idxPages_T_863_addr >= 6'h3e ? $random : idxPages[idxPages_T_863_addr];
  `endif
  assign idxPages_T_868_addr = 6'h3a;
  assign idxPages_T_868_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_868_data = idxPages[idxPages_T_868_addr];
  `else
  assign idxPages_T_868_data = idxPages_T_868_addr >= 6'h3e ? $random : idxPages[idxPages_T_868_addr];
  `endif
  assign idxPages_T_873_addr = 6'h3b;
  assign idxPages_T_873_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_873_data = idxPages[idxPages_T_873_addr];
  `else
  assign idxPages_T_873_data = idxPages_T_873_addr >= 6'h3e ? $random : idxPages[idxPages_T_873_addr];
  `endif
  assign idxPages_T_878_addr = 6'h3c;
  assign idxPages_T_878_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_878_data = idxPages[idxPages_T_878_addr];
  `else
  assign idxPages_T_878_data = idxPages_T_878_addr >= 6'h3e ? $random : idxPages[idxPages_T_878_addr];
  `endif
  assign idxPages_T_883_addr = 6'h3d;
  assign idxPages_T_883_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_883_data = idxPages[idxPages_T_883_addr];
  `else
  assign idxPages_T_883_data = idxPages_T_883_addr >= 6'h3e ? $random : idxPages[idxPages_T_883_addr];
  `endif
  assign idxPages_T_2874_data = idxPageUpdate;
  assign idxPages_T_2874_addr = T_2550;
  assign idxPages_T_2874_mask = r_btb_update_valid;
  assign idxPages_T_2874_en = r_btb_update_valid;
  assign tgts_T_3270_addr = {{5'd0}, 1'h0};
  assign tgts_T_3270_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3270_data = tgts[tgts_T_3270_addr];
  `else
  assign tgts_T_3270_data = tgts_T_3270_addr >= 6'h3e ? $random : tgts[tgts_T_3270_addr];
  `endif
  assign tgts_T_3272_addr = {{5'd0}, 1'h1};
  assign tgts_T_3272_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3272_data = tgts[tgts_T_3272_addr];
  `else
  assign tgts_T_3272_data = tgts_T_3272_addr >= 6'h3e ? $random : tgts[tgts_T_3272_addr];
  `endif
  assign tgts_T_3274_addr = {{4'd0}, 2'h2};
  assign tgts_T_3274_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3274_data = tgts[tgts_T_3274_addr];
  `else
  assign tgts_T_3274_data = tgts_T_3274_addr >= 6'h3e ? $random : tgts[tgts_T_3274_addr];
  `endif
  assign tgts_T_3276_addr = {{4'd0}, 2'h3};
  assign tgts_T_3276_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3276_data = tgts[tgts_T_3276_addr];
  `else
  assign tgts_T_3276_data = tgts_T_3276_addr >= 6'h3e ? $random : tgts[tgts_T_3276_addr];
  `endif
  assign tgts_T_3278_addr = {{3'd0}, 3'h4};
  assign tgts_T_3278_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3278_data = tgts[tgts_T_3278_addr];
  `else
  assign tgts_T_3278_data = tgts_T_3278_addr >= 6'h3e ? $random : tgts[tgts_T_3278_addr];
  `endif
  assign tgts_T_3280_addr = {{3'd0}, 3'h5};
  assign tgts_T_3280_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3280_data = tgts[tgts_T_3280_addr];
  `else
  assign tgts_T_3280_data = tgts_T_3280_addr >= 6'h3e ? $random : tgts[tgts_T_3280_addr];
  `endif
  assign tgts_T_3282_addr = {{3'd0}, 3'h6};
  assign tgts_T_3282_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3282_data = tgts[tgts_T_3282_addr];
  `else
  assign tgts_T_3282_data = tgts_T_3282_addr >= 6'h3e ? $random : tgts[tgts_T_3282_addr];
  `endif
  assign tgts_T_3284_addr = {{3'd0}, 3'h7};
  assign tgts_T_3284_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3284_data = tgts[tgts_T_3284_addr];
  `else
  assign tgts_T_3284_data = tgts_T_3284_addr >= 6'h3e ? $random : tgts[tgts_T_3284_addr];
  `endif
  assign tgts_T_3286_addr = {{2'd0}, 4'h8};
  assign tgts_T_3286_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3286_data = tgts[tgts_T_3286_addr];
  `else
  assign tgts_T_3286_data = tgts_T_3286_addr >= 6'h3e ? $random : tgts[tgts_T_3286_addr];
  `endif
  assign tgts_T_3288_addr = {{2'd0}, 4'h9};
  assign tgts_T_3288_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3288_data = tgts[tgts_T_3288_addr];
  `else
  assign tgts_T_3288_data = tgts_T_3288_addr >= 6'h3e ? $random : tgts[tgts_T_3288_addr];
  `endif
  assign tgts_T_3290_addr = {{2'd0}, 4'ha};
  assign tgts_T_3290_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3290_data = tgts[tgts_T_3290_addr];
  `else
  assign tgts_T_3290_data = tgts_T_3290_addr >= 6'h3e ? $random : tgts[tgts_T_3290_addr];
  `endif
  assign tgts_T_3292_addr = {{2'd0}, 4'hb};
  assign tgts_T_3292_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3292_data = tgts[tgts_T_3292_addr];
  `else
  assign tgts_T_3292_data = tgts_T_3292_addr >= 6'h3e ? $random : tgts[tgts_T_3292_addr];
  `endif
  assign tgts_T_3294_addr = {{2'd0}, 4'hc};
  assign tgts_T_3294_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3294_data = tgts[tgts_T_3294_addr];
  `else
  assign tgts_T_3294_data = tgts_T_3294_addr >= 6'h3e ? $random : tgts[tgts_T_3294_addr];
  `endif
  assign tgts_T_3296_addr = {{2'd0}, 4'hd};
  assign tgts_T_3296_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3296_data = tgts[tgts_T_3296_addr];
  `else
  assign tgts_T_3296_data = tgts_T_3296_addr >= 6'h3e ? $random : tgts[tgts_T_3296_addr];
  `endif
  assign tgts_T_3298_addr = {{2'd0}, 4'he};
  assign tgts_T_3298_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3298_data = tgts[tgts_T_3298_addr];
  `else
  assign tgts_T_3298_data = tgts_T_3298_addr >= 6'h3e ? $random : tgts[tgts_T_3298_addr];
  `endif
  assign tgts_T_3300_addr = {{2'd0}, 4'hf};
  assign tgts_T_3300_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3300_data = tgts[tgts_T_3300_addr];
  `else
  assign tgts_T_3300_data = tgts_T_3300_addr >= 6'h3e ? $random : tgts[tgts_T_3300_addr];
  `endif
  assign tgts_T_3302_addr = {{1'd0}, 5'h10};
  assign tgts_T_3302_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3302_data = tgts[tgts_T_3302_addr];
  `else
  assign tgts_T_3302_data = tgts_T_3302_addr >= 6'h3e ? $random : tgts[tgts_T_3302_addr];
  `endif
  assign tgts_T_3304_addr = {{1'd0}, 5'h11};
  assign tgts_T_3304_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3304_data = tgts[tgts_T_3304_addr];
  `else
  assign tgts_T_3304_data = tgts_T_3304_addr >= 6'h3e ? $random : tgts[tgts_T_3304_addr];
  `endif
  assign tgts_T_3306_addr = {{1'd0}, 5'h12};
  assign tgts_T_3306_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3306_data = tgts[tgts_T_3306_addr];
  `else
  assign tgts_T_3306_data = tgts_T_3306_addr >= 6'h3e ? $random : tgts[tgts_T_3306_addr];
  `endif
  assign tgts_T_3308_addr = {{1'd0}, 5'h13};
  assign tgts_T_3308_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3308_data = tgts[tgts_T_3308_addr];
  `else
  assign tgts_T_3308_data = tgts_T_3308_addr >= 6'h3e ? $random : tgts[tgts_T_3308_addr];
  `endif
  assign tgts_T_3310_addr = {{1'd0}, 5'h14};
  assign tgts_T_3310_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3310_data = tgts[tgts_T_3310_addr];
  `else
  assign tgts_T_3310_data = tgts_T_3310_addr >= 6'h3e ? $random : tgts[tgts_T_3310_addr];
  `endif
  assign tgts_T_3312_addr = {{1'd0}, 5'h15};
  assign tgts_T_3312_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3312_data = tgts[tgts_T_3312_addr];
  `else
  assign tgts_T_3312_data = tgts_T_3312_addr >= 6'h3e ? $random : tgts[tgts_T_3312_addr];
  `endif
  assign tgts_T_3314_addr = {{1'd0}, 5'h16};
  assign tgts_T_3314_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3314_data = tgts[tgts_T_3314_addr];
  `else
  assign tgts_T_3314_data = tgts_T_3314_addr >= 6'h3e ? $random : tgts[tgts_T_3314_addr];
  `endif
  assign tgts_T_3316_addr = {{1'd0}, 5'h17};
  assign tgts_T_3316_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3316_data = tgts[tgts_T_3316_addr];
  `else
  assign tgts_T_3316_data = tgts_T_3316_addr >= 6'h3e ? $random : tgts[tgts_T_3316_addr];
  `endif
  assign tgts_T_3318_addr = {{1'd0}, 5'h18};
  assign tgts_T_3318_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3318_data = tgts[tgts_T_3318_addr];
  `else
  assign tgts_T_3318_data = tgts_T_3318_addr >= 6'h3e ? $random : tgts[tgts_T_3318_addr];
  `endif
  assign tgts_T_3320_addr = {{1'd0}, 5'h19};
  assign tgts_T_3320_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3320_data = tgts[tgts_T_3320_addr];
  `else
  assign tgts_T_3320_data = tgts_T_3320_addr >= 6'h3e ? $random : tgts[tgts_T_3320_addr];
  `endif
  assign tgts_T_3322_addr = {{1'd0}, 5'h1a};
  assign tgts_T_3322_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3322_data = tgts[tgts_T_3322_addr];
  `else
  assign tgts_T_3322_data = tgts_T_3322_addr >= 6'h3e ? $random : tgts[tgts_T_3322_addr];
  `endif
  assign tgts_T_3324_addr = {{1'd0}, 5'h1b};
  assign tgts_T_3324_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3324_data = tgts[tgts_T_3324_addr];
  `else
  assign tgts_T_3324_data = tgts_T_3324_addr >= 6'h3e ? $random : tgts[tgts_T_3324_addr];
  `endif
  assign tgts_T_3326_addr = {{1'd0}, 5'h1c};
  assign tgts_T_3326_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3326_data = tgts[tgts_T_3326_addr];
  `else
  assign tgts_T_3326_data = tgts_T_3326_addr >= 6'h3e ? $random : tgts[tgts_T_3326_addr];
  `endif
  assign tgts_T_3328_addr = {{1'd0}, 5'h1d};
  assign tgts_T_3328_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3328_data = tgts[tgts_T_3328_addr];
  `else
  assign tgts_T_3328_data = tgts_T_3328_addr >= 6'h3e ? $random : tgts[tgts_T_3328_addr];
  `endif
  assign tgts_T_3330_addr = {{1'd0}, 5'h1e};
  assign tgts_T_3330_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3330_data = tgts[tgts_T_3330_addr];
  `else
  assign tgts_T_3330_data = tgts_T_3330_addr >= 6'h3e ? $random : tgts[tgts_T_3330_addr];
  `endif
  assign tgts_T_3332_addr = {{1'd0}, 5'h1f};
  assign tgts_T_3332_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3332_data = tgts[tgts_T_3332_addr];
  `else
  assign tgts_T_3332_data = tgts_T_3332_addr >= 6'h3e ? $random : tgts[tgts_T_3332_addr];
  `endif
  assign tgts_T_3334_addr = 6'h20;
  assign tgts_T_3334_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3334_data = tgts[tgts_T_3334_addr];
  `else
  assign tgts_T_3334_data = tgts_T_3334_addr >= 6'h3e ? $random : tgts[tgts_T_3334_addr];
  `endif
  assign tgts_T_3336_addr = 6'h21;
  assign tgts_T_3336_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3336_data = tgts[tgts_T_3336_addr];
  `else
  assign tgts_T_3336_data = tgts_T_3336_addr >= 6'h3e ? $random : tgts[tgts_T_3336_addr];
  `endif
  assign tgts_T_3338_addr = 6'h22;
  assign tgts_T_3338_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3338_data = tgts[tgts_T_3338_addr];
  `else
  assign tgts_T_3338_data = tgts_T_3338_addr >= 6'h3e ? $random : tgts[tgts_T_3338_addr];
  `endif
  assign tgts_T_3340_addr = 6'h23;
  assign tgts_T_3340_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3340_data = tgts[tgts_T_3340_addr];
  `else
  assign tgts_T_3340_data = tgts_T_3340_addr >= 6'h3e ? $random : tgts[tgts_T_3340_addr];
  `endif
  assign tgts_T_3342_addr = 6'h24;
  assign tgts_T_3342_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3342_data = tgts[tgts_T_3342_addr];
  `else
  assign tgts_T_3342_data = tgts_T_3342_addr >= 6'h3e ? $random : tgts[tgts_T_3342_addr];
  `endif
  assign tgts_T_3344_addr = 6'h25;
  assign tgts_T_3344_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3344_data = tgts[tgts_T_3344_addr];
  `else
  assign tgts_T_3344_data = tgts_T_3344_addr >= 6'h3e ? $random : tgts[tgts_T_3344_addr];
  `endif
  assign tgts_T_3346_addr = 6'h26;
  assign tgts_T_3346_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3346_data = tgts[tgts_T_3346_addr];
  `else
  assign tgts_T_3346_data = tgts_T_3346_addr >= 6'h3e ? $random : tgts[tgts_T_3346_addr];
  `endif
  assign tgts_T_3348_addr = 6'h27;
  assign tgts_T_3348_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3348_data = tgts[tgts_T_3348_addr];
  `else
  assign tgts_T_3348_data = tgts_T_3348_addr >= 6'h3e ? $random : tgts[tgts_T_3348_addr];
  `endif
  assign tgts_T_3350_addr = 6'h28;
  assign tgts_T_3350_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3350_data = tgts[tgts_T_3350_addr];
  `else
  assign tgts_T_3350_data = tgts_T_3350_addr >= 6'h3e ? $random : tgts[tgts_T_3350_addr];
  `endif
  assign tgts_T_3352_addr = 6'h29;
  assign tgts_T_3352_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3352_data = tgts[tgts_T_3352_addr];
  `else
  assign tgts_T_3352_data = tgts_T_3352_addr >= 6'h3e ? $random : tgts[tgts_T_3352_addr];
  `endif
  assign tgts_T_3354_addr = 6'h2a;
  assign tgts_T_3354_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3354_data = tgts[tgts_T_3354_addr];
  `else
  assign tgts_T_3354_data = tgts_T_3354_addr >= 6'h3e ? $random : tgts[tgts_T_3354_addr];
  `endif
  assign tgts_T_3356_addr = 6'h2b;
  assign tgts_T_3356_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3356_data = tgts[tgts_T_3356_addr];
  `else
  assign tgts_T_3356_data = tgts_T_3356_addr >= 6'h3e ? $random : tgts[tgts_T_3356_addr];
  `endif
  assign tgts_T_3358_addr = 6'h2c;
  assign tgts_T_3358_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3358_data = tgts[tgts_T_3358_addr];
  `else
  assign tgts_T_3358_data = tgts_T_3358_addr >= 6'h3e ? $random : tgts[tgts_T_3358_addr];
  `endif
  assign tgts_T_3360_addr = 6'h2d;
  assign tgts_T_3360_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3360_data = tgts[tgts_T_3360_addr];
  `else
  assign tgts_T_3360_data = tgts_T_3360_addr >= 6'h3e ? $random : tgts[tgts_T_3360_addr];
  `endif
  assign tgts_T_3362_addr = 6'h2e;
  assign tgts_T_3362_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3362_data = tgts[tgts_T_3362_addr];
  `else
  assign tgts_T_3362_data = tgts_T_3362_addr >= 6'h3e ? $random : tgts[tgts_T_3362_addr];
  `endif
  assign tgts_T_3364_addr = 6'h2f;
  assign tgts_T_3364_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3364_data = tgts[tgts_T_3364_addr];
  `else
  assign tgts_T_3364_data = tgts_T_3364_addr >= 6'h3e ? $random : tgts[tgts_T_3364_addr];
  `endif
  assign tgts_T_3366_addr = 6'h30;
  assign tgts_T_3366_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3366_data = tgts[tgts_T_3366_addr];
  `else
  assign tgts_T_3366_data = tgts_T_3366_addr >= 6'h3e ? $random : tgts[tgts_T_3366_addr];
  `endif
  assign tgts_T_3368_addr = 6'h31;
  assign tgts_T_3368_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3368_data = tgts[tgts_T_3368_addr];
  `else
  assign tgts_T_3368_data = tgts_T_3368_addr >= 6'h3e ? $random : tgts[tgts_T_3368_addr];
  `endif
  assign tgts_T_3370_addr = 6'h32;
  assign tgts_T_3370_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3370_data = tgts[tgts_T_3370_addr];
  `else
  assign tgts_T_3370_data = tgts_T_3370_addr >= 6'h3e ? $random : tgts[tgts_T_3370_addr];
  `endif
  assign tgts_T_3372_addr = 6'h33;
  assign tgts_T_3372_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3372_data = tgts[tgts_T_3372_addr];
  `else
  assign tgts_T_3372_data = tgts_T_3372_addr >= 6'h3e ? $random : tgts[tgts_T_3372_addr];
  `endif
  assign tgts_T_3374_addr = 6'h34;
  assign tgts_T_3374_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3374_data = tgts[tgts_T_3374_addr];
  `else
  assign tgts_T_3374_data = tgts_T_3374_addr >= 6'h3e ? $random : tgts[tgts_T_3374_addr];
  `endif
  assign tgts_T_3376_addr = 6'h35;
  assign tgts_T_3376_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3376_data = tgts[tgts_T_3376_addr];
  `else
  assign tgts_T_3376_data = tgts_T_3376_addr >= 6'h3e ? $random : tgts[tgts_T_3376_addr];
  `endif
  assign tgts_T_3378_addr = 6'h36;
  assign tgts_T_3378_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3378_data = tgts[tgts_T_3378_addr];
  `else
  assign tgts_T_3378_data = tgts_T_3378_addr >= 6'h3e ? $random : tgts[tgts_T_3378_addr];
  `endif
  assign tgts_T_3380_addr = 6'h37;
  assign tgts_T_3380_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3380_data = tgts[tgts_T_3380_addr];
  `else
  assign tgts_T_3380_data = tgts_T_3380_addr >= 6'h3e ? $random : tgts[tgts_T_3380_addr];
  `endif
  assign tgts_T_3382_addr = 6'h38;
  assign tgts_T_3382_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3382_data = tgts[tgts_T_3382_addr];
  `else
  assign tgts_T_3382_data = tgts_T_3382_addr >= 6'h3e ? $random : tgts[tgts_T_3382_addr];
  `endif
  assign tgts_T_3384_addr = 6'h39;
  assign tgts_T_3384_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3384_data = tgts[tgts_T_3384_addr];
  `else
  assign tgts_T_3384_data = tgts_T_3384_addr >= 6'h3e ? $random : tgts[tgts_T_3384_addr];
  `endif
  assign tgts_T_3386_addr = 6'h3a;
  assign tgts_T_3386_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3386_data = tgts[tgts_T_3386_addr];
  `else
  assign tgts_T_3386_data = tgts_T_3386_addr >= 6'h3e ? $random : tgts[tgts_T_3386_addr];
  `endif
  assign tgts_T_3388_addr = 6'h3b;
  assign tgts_T_3388_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3388_data = tgts[tgts_T_3388_addr];
  `else
  assign tgts_T_3388_data = tgts_T_3388_addr >= 6'h3e ? $random : tgts[tgts_T_3388_addr];
  `endif
  assign tgts_T_3390_addr = 6'h3c;
  assign tgts_T_3390_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3390_data = tgts[tgts_T_3390_addr];
  `else
  assign tgts_T_3390_data = tgts_T_3390_addr >= 6'h3e ? $random : tgts[tgts_T_3390_addr];
  `endif
  assign tgts_T_3392_addr = 6'h3d;
  assign tgts_T_3392_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3392_data = tgts[tgts_T_3392_addr];
  `else
  assign tgts_T_3392_data = tgts_T_3392_addr >= 6'h3e ? $random : tgts[tgts_T_3392_addr];
  `endif
  assign tgts_T_2873_data = io_req_bits_addr[11:0];
  assign tgts_T_2873_addr = T_2550;
  assign tgts_T_2873_mask = r_btb_update_valid;
  assign tgts_T_2873_en = r_btb_update_valid;
  assign tgtPages_T_888_addr = {{5'd0}, 1'h0};
  assign tgtPages_T_888_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_888_data = tgtPages[tgtPages_T_888_addr];
  `else
  assign tgtPages_T_888_data = tgtPages_T_888_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_888_addr];
  `endif
  assign tgtPages_T_893_addr = {{5'd0}, 1'h1};
  assign tgtPages_T_893_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_893_data = tgtPages[tgtPages_T_893_addr];
  `else
  assign tgtPages_T_893_data = tgtPages_T_893_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_893_addr];
  `endif
  assign tgtPages_T_898_addr = {{4'd0}, 2'h2};
  assign tgtPages_T_898_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_898_data = tgtPages[tgtPages_T_898_addr];
  `else
  assign tgtPages_T_898_data = tgtPages_T_898_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_898_addr];
  `endif
  assign tgtPages_T_903_addr = {{4'd0}, 2'h3};
  assign tgtPages_T_903_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_903_data = tgtPages[tgtPages_T_903_addr];
  `else
  assign tgtPages_T_903_data = tgtPages_T_903_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_903_addr];
  `endif
  assign tgtPages_T_908_addr = {{3'd0}, 3'h4};
  assign tgtPages_T_908_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_908_data = tgtPages[tgtPages_T_908_addr];
  `else
  assign tgtPages_T_908_data = tgtPages_T_908_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_908_addr];
  `endif
  assign tgtPages_T_913_addr = {{3'd0}, 3'h5};
  assign tgtPages_T_913_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_913_data = tgtPages[tgtPages_T_913_addr];
  `else
  assign tgtPages_T_913_data = tgtPages_T_913_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_913_addr];
  `endif
  assign tgtPages_T_918_addr = {{3'd0}, 3'h6};
  assign tgtPages_T_918_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_918_data = tgtPages[tgtPages_T_918_addr];
  `else
  assign tgtPages_T_918_data = tgtPages_T_918_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_918_addr];
  `endif
  assign tgtPages_T_923_addr = {{3'd0}, 3'h7};
  assign tgtPages_T_923_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_923_data = tgtPages[tgtPages_T_923_addr];
  `else
  assign tgtPages_T_923_data = tgtPages_T_923_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_923_addr];
  `endif
  assign tgtPages_T_928_addr = {{2'd0}, 4'h8};
  assign tgtPages_T_928_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_928_data = tgtPages[tgtPages_T_928_addr];
  `else
  assign tgtPages_T_928_data = tgtPages_T_928_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_928_addr];
  `endif
  assign tgtPages_T_933_addr = {{2'd0}, 4'h9};
  assign tgtPages_T_933_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_933_data = tgtPages[tgtPages_T_933_addr];
  `else
  assign tgtPages_T_933_data = tgtPages_T_933_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_933_addr];
  `endif
  assign tgtPages_T_938_addr = {{2'd0}, 4'ha};
  assign tgtPages_T_938_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_938_data = tgtPages[tgtPages_T_938_addr];
  `else
  assign tgtPages_T_938_data = tgtPages_T_938_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_938_addr];
  `endif
  assign tgtPages_T_943_addr = {{2'd0}, 4'hb};
  assign tgtPages_T_943_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_943_data = tgtPages[tgtPages_T_943_addr];
  `else
  assign tgtPages_T_943_data = tgtPages_T_943_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_943_addr];
  `endif
  assign tgtPages_T_948_addr = {{2'd0}, 4'hc};
  assign tgtPages_T_948_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_948_data = tgtPages[tgtPages_T_948_addr];
  `else
  assign tgtPages_T_948_data = tgtPages_T_948_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_948_addr];
  `endif
  assign tgtPages_T_953_addr = {{2'd0}, 4'hd};
  assign tgtPages_T_953_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_953_data = tgtPages[tgtPages_T_953_addr];
  `else
  assign tgtPages_T_953_data = tgtPages_T_953_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_953_addr];
  `endif
  assign tgtPages_T_958_addr = {{2'd0}, 4'he};
  assign tgtPages_T_958_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_958_data = tgtPages[tgtPages_T_958_addr];
  `else
  assign tgtPages_T_958_data = tgtPages_T_958_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_958_addr];
  `endif
  assign tgtPages_T_963_addr = {{2'd0}, 4'hf};
  assign tgtPages_T_963_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_963_data = tgtPages[tgtPages_T_963_addr];
  `else
  assign tgtPages_T_963_data = tgtPages_T_963_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_963_addr];
  `endif
  assign tgtPages_T_968_addr = {{1'd0}, 5'h10};
  assign tgtPages_T_968_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_968_data = tgtPages[tgtPages_T_968_addr];
  `else
  assign tgtPages_T_968_data = tgtPages_T_968_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_968_addr];
  `endif
  assign tgtPages_T_973_addr = {{1'd0}, 5'h11};
  assign tgtPages_T_973_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_973_data = tgtPages[tgtPages_T_973_addr];
  `else
  assign tgtPages_T_973_data = tgtPages_T_973_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_973_addr];
  `endif
  assign tgtPages_T_978_addr = {{1'd0}, 5'h12};
  assign tgtPages_T_978_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_978_data = tgtPages[tgtPages_T_978_addr];
  `else
  assign tgtPages_T_978_data = tgtPages_T_978_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_978_addr];
  `endif
  assign tgtPages_T_983_addr = {{1'd0}, 5'h13};
  assign tgtPages_T_983_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_983_data = tgtPages[tgtPages_T_983_addr];
  `else
  assign tgtPages_T_983_data = tgtPages_T_983_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_983_addr];
  `endif
  assign tgtPages_T_988_addr = {{1'd0}, 5'h14};
  assign tgtPages_T_988_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_988_data = tgtPages[tgtPages_T_988_addr];
  `else
  assign tgtPages_T_988_data = tgtPages_T_988_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_988_addr];
  `endif
  assign tgtPages_T_993_addr = {{1'd0}, 5'h15};
  assign tgtPages_T_993_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_993_data = tgtPages[tgtPages_T_993_addr];
  `else
  assign tgtPages_T_993_data = tgtPages_T_993_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_993_addr];
  `endif
  assign tgtPages_T_998_addr = {{1'd0}, 5'h16};
  assign tgtPages_T_998_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_998_data = tgtPages[tgtPages_T_998_addr];
  `else
  assign tgtPages_T_998_data = tgtPages_T_998_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_998_addr];
  `endif
  assign tgtPages_T_1003_addr = {{1'd0}, 5'h17};
  assign tgtPages_T_1003_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1003_data = tgtPages[tgtPages_T_1003_addr];
  `else
  assign tgtPages_T_1003_data = tgtPages_T_1003_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1003_addr];
  `endif
  assign tgtPages_T_1008_addr = {{1'd0}, 5'h18};
  assign tgtPages_T_1008_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1008_data = tgtPages[tgtPages_T_1008_addr];
  `else
  assign tgtPages_T_1008_data = tgtPages_T_1008_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1008_addr];
  `endif
  assign tgtPages_T_1013_addr = {{1'd0}, 5'h19};
  assign tgtPages_T_1013_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1013_data = tgtPages[tgtPages_T_1013_addr];
  `else
  assign tgtPages_T_1013_data = tgtPages_T_1013_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1013_addr];
  `endif
  assign tgtPages_T_1018_addr = {{1'd0}, 5'h1a};
  assign tgtPages_T_1018_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1018_data = tgtPages[tgtPages_T_1018_addr];
  `else
  assign tgtPages_T_1018_data = tgtPages_T_1018_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1018_addr];
  `endif
  assign tgtPages_T_1023_addr = {{1'd0}, 5'h1b};
  assign tgtPages_T_1023_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1023_data = tgtPages[tgtPages_T_1023_addr];
  `else
  assign tgtPages_T_1023_data = tgtPages_T_1023_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1023_addr];
  `endif
  assign tgtPages_T_1028_addr = {{1'd0}, 5'h1c};
  assign tgtPages_T_1028_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1028_data = tgtPages[tgtPages_T_1028_addr];
  `else
  assign tgtPages_T_1028_data = tgtPages_T_1028_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1028_addr];
  `endif
  assign tgtPages_T_1033_addr = {{1'd0}, 5'h1d};
  assign tgtPages_T_1033_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1033_data = tgtPages[tgtPages_T_1033_addr];
  `else
  assign tgtPages_T_1033_data = tgtPages_T_1033_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1033_addr];
  `endif
  assign tgtPages_T_1038_addr = {{1'd0}, 5'h1e};
  assign tgtPages_T_1038_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1038_data = tgtPages[tgtPages_T_1038_addr];
  `else
  assign tgtPages_T_1038_data = tgtPages_T_1038_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1038_addr];
  `endif
  assign tgtPages_T_1043_addr = {{1'd0}, 5'h1f};
  assign tgtPages_T_1043_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1043_data = tgtPages[tgtPages_T_1043_addr];
  `else
  assign tgtPages_T_1043_data = tgtPages_T_1043_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1043_addr];
  `endif
  assign tgtPages_T_1048_addr = 6'h20;
  assign tgtPages_T_1048_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1048_data = tgtPages[tgtPages_T_1048_addr];
  `else
  assign tgtPages_T_1048_data = tgtPages_T_1048_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1048_addr];
  `endif
  assign tgtPages_T_1053_addr = 6'h21;
  assign tgtPages_T_1053_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1053_data = tgtPages[tgtPages_T_1053_addr];
  `else
  assign tgtPages_T_1053_data = tgtPages_T_1053_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1053_addr];
  `endif
  assign tgtPages_T_1058_addr = 6'h22;
  assign tgtPages_T_1058_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1058_data = tgtPages[tgtPages_T_1058_addr];
  `else
  assign tgtPages_T_1058_data = tgtPages_T_1058_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1058_addr];
  `endif
  assign tgtPages_T_1063_addr = 6'h23;
  assign tgtPages_T_1063_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1063_data = tgtPages[tgtPages_T_1063_addr];
  `else
  assign tgtPages_T_1063_data = tgtPages_T_1063_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1063_addr];
  `endif
  assign tgtPages_T_1068_addr = 6'h24;
  assign tgtPages_T_1068_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1068_data = tgtPages[tgtPages_T_1068_addr];
  `else
  assign tgtPages_T_1068_data = tgtPages_T_1068_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1068_addr];
  `endif
  assign tgtPages_T_1073_addr = 6'h25;
  assign tgtPages_T_1073_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1073_data = tgtPages[tgtPages_T_1073_addr];
  `else
  assign tgtPages_T_1073_data = tgtPages_T_1073_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1073_addr];
  `endif
  assign tgtPages_T_1078_addr = 6'h26;
  assign tgtPages_T_1078_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1078_data = tgtPages[tgtPages_T_1078_addr];
  `else
  assign tgtPages_T_1078_data = tgtPages_T_1078_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1078_addr];
  `endif
  assign tgtPages_T_1083_addr = 6'h27;
  assign tgtPages_T_1083_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1083_data = tgtPages[tgtPages_T_1083_addr];
  `else
  assign tgtPages_T_1083_data = tgtPages_T_1083_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1083_addr];
  `endif
  assign tgtPages_T_1088_addr = 6'h28;
  assign tgtPages_T_1088_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1088_data = tgtPages[tgtPages_T_1088_addr];
  `else
  assign tgtPages_T_1088_data = tgtPages_T_1088_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1088_addr];
  `endif
  assign tgtPages_T_1093_addr = 6'h29;
  assign tgtPages_T_1093_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1093_data = tgtPages[tgtPages_T_1093_addr];
  `else
  assign tgtPages_T_1093_data = tgtPages_T_1093_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1093_addr];
  `endif
  assign tgtPages_T_1098_addr = 6'h2a;
  assign tgtPages_T_1098_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1098_data = tgtPages[tgtPages_T_1098_addr];
  `else
  assign tgtPages_T_1098_data = tgtPages_T_1098_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1098_addr];
  `endif
  assign tgtPages_T_1103_addr = 6'h2b;
  assign tgtPages_T_1103_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1103_data = tgtPages[tgtPages_T_1103_addr];
  `else
  assign tgtPages_T_1103_data = tgtPages_T_1103_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1103_addr];
  `endif
  assign tgtPages_T_1108_addr = 6'h2c;
  assign tgtPages_T_1108_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1108_data = tgtPages[tgtPages_T_1108_addr];
  `else
  assign tgtPages_T_1108_data = tgtPages_T_1108_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1108_addr];
  `endif
  assign tgtPages_T_1113_addr = 6'h2d;
  assign tgtPages_T_1113_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1113_data = tgtPages[tgtPages_T_1113_addr];
  `else
  assign tgtPages_T_1113_data = tgtPages_T_1113_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1113_addr];
  `endif
  assign tgtPages_T_1118_addr = 6'h2e;
  assign tgtPages_T_1118_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1118_data = tgtPages[tgtPages_T_1118_addr];
  `else
  assign tgtPages_T_1118_data = tgtPages_T_1118_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1118_addr];
  `endif
  assign tgtPages_T_1123_addr = 6'h2f;
  assign tgtPages_T_1123_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1123_data = tgtPages[tgtPages_T_1123_addr];
  `else
  assign tgtPages_T_1123_data = tgtPages_T_1123_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1123_addr];
  `endif
  assign tgtPages_T_1128_addr = 6'h30;
  assign tgtPages_T_1128_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1128_data = tgtPages[tgtPages_T_1128_addr];
  `else
  assign tgtPages_T_1128_data = tgtPages_T_1128_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1128_addr];
  `endif
  assign tgtPages_T_1133_addr = 6'h31;
  assign tgtPages_T_1133_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1133_data = tgtPages[tgtPages_T_1133_addr];
  `else
  assign tgtPages_T_1133_data = tgtPages_T_1133_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1133_addr];
  `endif
  assign tgtPages_T_1138_addr = 6'h32;
  assign tgtPages_T_1138_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1138_data = tgtPages[tgtPages_T_1138_addr];
  `else
  assign tgtPages_T_1138_data = tgtPages_T_1138_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1138_addr];
  `endif
  assign tgtPages_T_1143_addr = 6'h33;
  assign tgtPages_T_1143_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1143_data = tgtPages[tgtPages_T_1143_addr];
  `else
  assign tgtPages_T_1143_data = tgtPages_T_1143_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1143_addr];
  `endif
  assign tgtPages_T_1148_addr = 6'h34;
  assign tgtPages_T_1148_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1148_data = tgtPages[tgtPages_T_1148_addr];
  `else
  assign tgtPages_T_1148_data = tgtPages_T_1148_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1148_addr];
  `endif
  assign tgtPages_T_1153_addr = 6'h35;
  assign tgtPages_T_1153_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1153_data = tgtPages[tgtPages_T_1153_addr];
  `else
  assign tgtPages_T_1153_data = tgtPages_T_1153_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1153_addr];
  `endif
  assign tgtPages_T_1158_addr = 6'h36;
  assign tgtPages_T_1158_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1158_data = tgtPages[tgtPages_T_1158_addr];
  `else
  assign tgtPages_T_1158_data = tgtPages_T_1158_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1158_addr];
  `endif
  assign tgtPages_T_1163_addr = 6'h37;
  assign tgtPages_T_1163_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1163_data = tgtPages[tgtPages_T_1163_addr];
  `else
  assign tgtPages_T_1163_data = tgtPages_T_1163_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1163_addr];
  `endif
  assign tgtPages_T_1168_addr = 6'h38;
  assign tgtPages_T_1168_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1168_data = tgtPages[tgtPages_T_1168_addr];
  `else
  assign tgtPages_T_1168_data = tgtPages_T_1168_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1168_addr];
  `endif
  assign tgtPages_T_1173_addr = 6'h39;
  assign tgtPages_T_1173_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1173_data = tgtPages[tgtPages_T_1173_addr];
  `else
  assign tgtPages_T_1173_data = tgtPages_T_1173_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1173_addr];
  `endif
  assign tgtPages_T_1178_addr = 6'h3a;
  assign tgtPages_T_1178_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1178_data = tgtPages[tgtPages_T_1178_addr];
  `else
  assign tgtPages_T_1178_data = tgtPages_T_1178_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1178_addr];
  `endif
  assign tgtPages_T_1183_addr = 6'h3b;
  assign tgtPages_T_1183_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1183_data = tgtPages[tgtPages_T_1183_addr];
  `else
  assign tgtPages_T_1183_data = tgtPages_T_1183_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1183_addr];
  `endif
  assign tgtPages_T_1188_addr = 6'h3c;
  assign tgtPages_T_1188_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1188_data = tgtPages[tgtPages_T_1188_addr];
  `else
  assign tgtPages_T_1188_data = tgtPages_T_1188_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1188_addr];
  `endif
  assign tgtPages_T_1193_addr = 6'h3d;
  assign tgtPages_T_1193_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1193_data = tgtPages[tgtPages_T_1193_addr];
  `else
  assign tgtPages_T_1193_data = tgtPages_T_1193_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1193_addr];
  `endif
  assign tgtPages_T_2875_data = tgtPageUpdate;
  assign tgtPages_T_2875_addr = T_2550;
  assign tgtPages_T_2875_mask = r_btb_update_valid;
  assign tgtPages_T_2875_en = r_btb_update_valid;
  assign pages_T_1400_addr = {{2'd0}, 1'h0};
  assign pages_T_1400_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1400_data = pages[pages_T_1400_addr];
  `else
  assign pages_T_1400_data = pages_T_1400_addr >= 3'h6 ? $random : pages[pages_T_1400_addr];
  `endif
  assign pages_T_1403_addr = {{2'd0}, 1'h1};
  assign pages_T_1403_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1403_data = pages[pages_T_1403_addr];
  `else
  assign pages_T_1403_data = pages_T_1403_addr >= 3'h6 ? $random : pages[pages_T_1403_addr];
  `endif
  assign pages_T_1406_addr = {{1'd0}, 2'h2};
  assign pages_T_1406_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1406_data = pages[pages_T_1406_addr];
  `else
  assign pages_T_1406_data = pages_T_1406_addr >= 3'h6 ? $random : pages[pages_T_1406_addr];
  `endif
  assign pages_T_1409_addr = {{1'd0}, 2'h3};
  assign pages_T_1409_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1409_data = pages[pages_T_1409_addr];
  `else
  assign pages_T_1409_data = pages_T_1409_addr >= 3'h6 ? $random : pages[pages_T_1409_addr];
  `endif
  assign pages_T_1412_addr = 3'h4;
  assign pages_T_1412_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1412_data = pages[pages_T_1412_addr];
  `else
  assign pages_T_1412_data = pages_T_1412_addr >= 3'h6 ? $random : pages[pages_T_1412_addr];
  `endif
  assign pages_T_1415_addr = 3'h5;
  assign pages_T_1415_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1415_data = pages[pages_T_1415_addr];
  `else
  assign pages_T_1415_data = pages_T_1415_addr >= 3'h6 ? $random : pages[pages_T_1415_addr];
  `endif
  assign pages_T_1941_addr = {{2'd0}, 1'h0};
  assign pages_T_1941_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1941_data = pages[pages_T_1941_addr];
  `else
  assign pages_T_1941_data = pages_T_1941_addr >= 3'h6 ? $random : pages[pages_T_1941_addr];
  `endif
  assign pages_T_1944_addr = {{2'd0}, 1'h1};
  assign pages_T_1944_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1944_data = pages[pages_T_1944_addr];
  `else
  assign pages_T_1944_data = pages_T_1944_addr >= 3'h6 ? $random : pages[pages_T_1944_addr];
  `endif
  assign pages_T_1947_addr = {{1'd0}, 2'h2};
  assign pages_T_1947_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1947_data = pages[pages_T_1947_addr];
  `else
  assign pages_T_1947_data = pages_T_1947_addr >= 3'h6 ? $random : pages[pages_T_1947_addr];
  `endif
  assign pages_T_1950_addr = {{1'd0}, 2'h3};
  assign pages_T_1950_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1950_data = pages[pages_T_1950_addr];
  `else
  assign pages_T_1950_data = pages_T_1950_addr >= 3'h6 ? $random : pages[pages_T_1950_addr];
  `endif
  assign pages_T_1953_addr = 3'h4;
  assign pages_T_1953_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1953_data = pages[pages_T_1953_addr];
  `else
  assign pages_T_1953_data = pages_T_1953_addr >= 3'h6 ? $random : pages[pages_T_1953_addr];
  `endif
  assign pages_T_1956_addr = 3'h5;
  assign pages_T_1956_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1956_data = pages[pages_T_1956_addr];
  `else
  assign pages_T_1956_data = pages_T_1956_addr >= 3'h6 ? $random : pages[pages_T_1956_addr];
  `endif
  assign pages_T_3177_addr = {{2'd0}, 1'h0};
  assign pages_T_3177_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3177_data = pages[pages_T_3177_addr];
  `else
  assign pages_T_3177_data = pages_T_3177_addr >= 3'h6 ? $random : pages[pages_T_3177_addr];
  `endif
  assign pages_T_3179_addr = {{2'd0}, 1'h1};
  assign pages_T_3179_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3179_data = pages[pages_T_3179_addr];
  `else
  assign pages_T_3179_data = pages_T_3179_addr >= 3'h6 ? $random : pages[pages_T_3179_addr];
  `endif
  assign pages_T_3181_addr = {{1'd0}, 2'h2};
  assign pages_T_3181_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3181_data = pages[pages_T_3181_addr];
  `else
  assign pages_T_3181_data = pages_T_3181_addr >= 3'h6 ? $random : pages[pages_T_3181_addr];
  `endif
  assign pages_T_3183_addr = {{1'd0}, 2'h3};
  assign pages_T_3183_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3183_data = pages[pages_T_3183_addr];
  `else
  assign pages_T_3183_data = pages_T_3183_addr >= 3'h6 ? $random : pages[pages_T_3183_addr];
  `endif
  assign pages_T_3185_addr = 3'h4;
  assign pages_T_3185_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3185_data = pages[pages_T_3185_addr];
  `else
  assign pages_T_3185_data = pages_T_3185_addr >= 3'h6 ? $random : pages[pages_T_3185_addr];
  `endif
  assign pages_T_3187_addr = 3'h5;
  assign pages_T_3187_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3187_data = pages[pages_T_3187_addr];
  `else
  assign pages_T_3187_data = pages_T_3187_addr >= 3'h6 ? $random : pages[pages_T_3187_addr];
  `endif
  assign pages_T_2891_data = T_2887;
  assign pages_T_2891_addr = {{2'd0}, 1'h0};
  assign pages_T_2891_mask = GEN_393;
  assign pages_T_2891_en = GEN_393;
  assign pages_T_2895_data = T_2887;
  assign pages_T_2895_addr = {{1'd0}, 2'h2};
  assign pages_T_2895_mask = GEN_398;
  assign pages_T_2895_en = GEN_398;
  assign pages_T_2899_data = T_2887;
  assign pages_T_2899_addr = 3'h4;
  assign pages_T_2899_mask = GEN_403;
  assign pages_T_2899_en = GEN_403;
  assign pages_T_2907_data = T_2903;
  assign pages_T_2907_addr = {{2'd0}, 1'h1};
  assign pages_T_2907_mask = GEN_408;
  assign pages_T_2907_en = GEN_408;
  assign pages_T_2911_data = T_2903;
  assign pages_T_2911_addr = {{1'd0}, 2'h3};
  assign pages_T_2911_mask = GEN_413;
  assign pages_T_2911_en = GEN_413;
  assign pages_T_2915_data = T_2903;
  assign pages_T_2915_addr = 3'h5;
  assign pages_T_2915_mask = GEN_418;
  assign pages_T_2915_en = GEN_418;
  assign GEN_457 = {{7'd0}, 1'h1};
  assign T_580 = GEN_457 << idxPages_T_578_data;
  assign T_581 = T_580[5:0];
  assign T_585 = GEN_457 << idxPages_T_583_data;
  assign T_586 = T_585[5:0];
  assign T_590 = GEN_457 << idxPages_T_588_data;
  assign T_591 = T_590[5:0];
  assign T_595 = GEN_457 << idxPages_T_593_data;
  assign T_596 = T_595[5:0];
  assign T_600 = GEN_457 << idxPages_T_598_data;
  assign T_601 = T_600[5:0];
  assign T_605 = GEN_457 << idxPages_T_603_data;
  assign T_606 = T_605[5:0];
  assign T_610 = GEN_457 << idxPages_T_608_data;
  assign T_611 = T_610[5:0];
  assign T_615 = GEN_457 << idxPages_T_613_data;
  assign T_616 = T_615[5:0];
  assign T_620 = GEN_457 << idxPages_T_618_data;
  assign T_621 = T_620[5:0];
  assign T_625 = GEN_457 << idxPages_T_623_data;
  assign T_626 = T_625[5:0];
  assign T_630 = GEN_457 << idxPages_T_628_data;
  assign T_631 = T_630[5:0];
  assign T_635 = GEN_457 << idxPages_T_633_data;
  assign T_636 = T_635[5:0];
  assign T_640 = GEN_457 << idxPages_T_638_data;
  assign T_641 = T_640[5:0];
  assign T_645 = GEN_457 << idxPages_T_643_data;
  assign T_646 = T_645[5:0];
  assign T_650 = GEN_457 << idxPages_T_648_data;
  assign T_651 = T_650[5:0];
  assign T_655 = GEN_457 << idxPages_T_653_data;
  assign T_656 = T_655[5:0];
  assign T_660 = GEN_457 << idxPages_T_658_data;
  assign T_661 = T_660[5:0];
  assign T_665 = GEN_457 << idxPages_T_663_data;
  assign T_666 = T_665[5:0];
  assign T_670 = GEN_457 << idxPages_T_668_data;
  assign T_671 = T_670[5:0];
  assign T_675 = GEN_457 << idxPages_T_673_data;
  assign T_676 = T_675[5:0];
  assign T_680 = GEN_457 << idxPages_T_678_data;
  assign T_681 = T_680[5:0];
  assign T_685 = GEN_457 << idxPages_T_683_data;
  assign T_686 = T_685[5:0];
  assign T_690 = GEN_457 << idxPages_T_688_data;
  assign T_691 = T_690[5:0];
  assign T_695 = GEN_457 << idxPages_T_693_data;
  assign T_696 = T_695[5:0];
  assign T_700 = GEN_457 << idxPages_T_698_data;
  assign T_701 = T_700[5:0];
  assign T_705 = GEN_457 << idxPages_T_703_data;
  assign T_706 = T_705[5:0];
  assign T_710 = GEN_457 << idxPages_T_708_data;
  assign T_711 = T_710[5:0];
  assign T_715 = GEN_457 << idxPages_T_713_data;
  assign T_716 = T_715[5:0];
  assign T_720 = GEN_457 << idxPages_T_718_data;
  assign T_721 = T_720[5:0];
  assign T_725 = GEN_457 << idxPages_T_723_data;
  assign T_726 = T_725[5:0];
  assign T_730 = GEN_457 << idxPages_T_728_data;
  assign T_731 = T_730[5:0];
  assign T_735 = GEN_457 << idxPages_T_733_data;
  assign T_736 = T_735[5:0];
  assign T_740 = GEN_457 << idxPages_T_738_data;
  assign T_741 = T_740[5:0];
  assign T_745 = GEN_457 << idxPages_T_743_data;
  assign T_746 = T_745[5:0];
  assign T_750 = GEN_457 << idxPages_T_748_data;
  assign T_751 = T_750[5:0];
  assign T_755 = GEN_457 << idxPages_T_753_data;
  assign T_756 = T_755[5:0];
  assign T_760 = GEN_457 << idxPages_T_758_data;
  assign T_761 = T_760[5:0];
  assign T_765 = GEN_457 << idxPages_T_763_data;
  assign T_766 = T_765[5:0];
  assign T_770 = GEN_457 << idxPages_T_768_data;
  assign T_771 = T_770[5:0];
  assign T_775 = GEN_457 << idxPages_T_773_data;
  assign T_776 = T_775[5:0];
  assign T_780 = GEN_457 << idxPages_T_778_data;
  assign T_781 = T_780[5:0];
  assign T_785 = GEN_457 << idxPages_T_783_data;
  assign T_786 = T_785[5:0];
  assign T_790 = GEN_457 << idxPages_T_788_data;
  assign T_791 = T_790[5:0];
  assign T_795 = GEN_457 << idxPages_T_793_data;
  assign T_796 = T_795[5:0];
  assign T_800 = GEN_457 << idxPages_T_798_data;
  assign T_801 = T_800[5:0];
  assign T_805 = GEN_457 << idxPages_T_803_data;
  assign T_806 = T_805[5:0];
  assign T_810 = GEN_457 << idxPages_T_808_data;
  assign T_811 = T_810[5:0];
  assign T_815 = GEN_457 << idxPages_T_813_data;
  assign T_816 = T_815[5:0];
  assign T_820 = GEN_457 << idxPages_T_818_data;
  assign T_821 = T_820[5:0];
  assign T_825 = GEN_457 << idxPages_T_823_data;
  assign T_826 = T_825[5:0];
  assign T_830 = GEN_457 << idxPages_T_828_data;
  assign T_831 = T_830[5:0];
  assign T_835 = GEN_457 << idxPages_T_833_data;
  assign T_836 = T_835[5:0];
  assign T_840 = GEN_457 << idxPages_T_838_data;
  assign T_841 = T_840[5:0];
  assign T_845 = GEN_457 << idxPages_T_843_data;
  assign T_846 = T_845[5:0];
  assign T_850 = GEN_457 << idxPages_T_848_data;
  assign T_851 = T_850[5:0];
  assign T_855 = GEN_457 << idxPages_T_853_data;
  assign T_856 = T_855[5:0];
  assign T_860 = GEN_457 << idxPages_T_858_data;
  assign T_861 = T_860[5:0];
  assign T_865 = GEN_457 << idxPages_T_863_data;
  assign T_866 = T_865[5:0];
  assign T_870 = GEN_457 << idxPages_T_868_data;
  assign T_871 = T_870[5:0];
  assign T_875 = GEN_457 << idxPages_T_873_data;
  assign T_876 = T_875[5:0];
  assign T_880 = GEN_457 << idxPages_T_878_data;
  assign T_881 = T_880[5:0];
  assign T_885 = GEN_457 << idxPages_T_883_data;
  assign T_886 = T_885[5:0];
  assign T_890 = GEN_457 << tgtPages_T_888_data;
  assign T_891 = T_890[5:0];
  assign T_895 = GEN_457 << tgtPages_T_893_data;
  assign T_896 = T_895[5:0];
  assign T_900 = GEN_457 << tgtPages_T_898_data;
  assign T_901 = T_900[5:0];
  assign T_905 = GEN_457 << tgtPages_T_903_data;
  assign T_906 = T_905[5:0];
  assign T_910 = GEN_457 << tgtPages_T_908_data;
  assign T_911 = T_910[5:0];
  assign T_915 = GEN_457 << tgtPages_T_913_data;
  assign T_916 = T_915[5:0];
  assign T_920 = GEN_457 << tgtPages_T_918_data;
  assign T_921 = T_920[5:0];
  assign T_925 = GEN_457 << tgtPages_T_923_data;
  assign T_926 = T_925[5:0];
  assign T_930 = GEN_457 << tgtPages_T_928_data;
  assign T_931 = T_930[5:0];
  assign T_935 = GEN_457 << tgtPages_T_933_data;
  assign T_936 = T_935[5:0];
  assign T_940 = GEN_457 << tgtPages_T_938_data;
  assign T_941 = T_940[5:0];
  assign T_945 = GEN_457 << tgtPages_T_943_data;
  assign T_946 = T_945[5:0];
  assign T_950 = GEN_457 << tgtPages_T_948_data;
  assign T_951 = T_950[5:0];
  assign T_955 = GEN_457 << tgtPages_T_953_data;
  assign T_956 = T_955[5:0];
  assign T_960 = GEN_457 << tgtPages_T_958_data;
  assign T_961 = T_960[5:0];
  assign T_965 = GEN_457 << tgtPages_T_963_data;
  assign T_966 = T_965[5:0];
  assign T_970 = GEN_457 << tgtPages_T_968_data;
  assign T_971 = T_970[5:0];
  assign T_975 = GEN_457 << tgtPages_T_973_data;
  assign T_976 = T_975[5:0];
  assign T_980 = GEN_457 << tgtPages_T_978_data;
  assign T_981 = T_980[5:0];
  assign T_985 = GEN_457 << tgtPages_T_983_data;
  assign T_986 = T_985[5:0];
  assign T_990 = GEN_457 << tgtPages_T_988_data;
  assign T_991 = T_990[5:0];
  assign T_995 = GEN_457 << tgtPages_T_993_data;
  assign T_996 = T_995[5:0];
  assign T_1000 = GEN_457 << tgtPages_T_998_data;
  assign T_1001 = T_1000[5:0];
  assign T_1005 = GEN_457 << tgtPages_T_1003_data;
  assign T_1006 = T_1005[5:0];
  assign T_1010 = GEN_457 << tgtPages_T_1008_data;
  assign T_1011 = T_1010[5:0];
  assign T_1015 = GEN_457 << tgtPages_T_1013_data;
  assign T_1016 = T_1015[5:0];
  assign T_1020 = GEN_457 << tgtPages_T_1018_data;
  assign T_1021 = T_1020[5:0];
  assign T_1025 = GEN_457 << tgtPages_T_1023_data;
  assign T_1026 = T_1025[5:0];
  assign T_1030 = GEN_457 << tgtPages_T_1028_data;
  assign T_1031 = T_1030[5:0];
  assign T_1035 = GEN_457 << tgtPages_T_1033_data;
  assign T_1036 = T_1035[5:0];
  assign T_1040 = GEN_457 << tgtPages_T_1038_data;
  assign T_1041 = T_1040[5:0];
  assign T_1045 = GEN_457 << tgtPages_T_1043_data;
  assign T_1046 = T_1045[5:0];
  assign T_1050 = GEN_457 << tgtPages_T_1048_data;
  assign T_1051 = T_1050[5:0];
  assign T_1055 = GEN_457 << tgtPages_T_1053_data;
  assign T_1056 = T_1055[5:0];
  assign T_1060 = GEN_457 << tgtPages_T_1058_data;
  assign T_1061 = T_1060[5:0];
  assign T_1065 = GEN_457 << tgtPages_T_1063_data;
  assign T_1066 = T_1065[5:0];
  assign T_1070 = GEN_457 << tgtPages_T_1068_data;
  assign T_1071 = T_1070[5:0];
  assign T_1075 = GEN_457 << tgtPages_T_1073_data;
  assign T_1076 = T_1075[5:0];
  assign T_1080 = GEN_457 << tgtPages_T_1078_data;
  assign T_1081 = T_1080[5:0];
  assign T_1085 = GEN_457 << tgtPages_T_1083_data;
  assign T_1086 = T_1085[5:0];
  assign T_1090 = GEN_457 << tgtPages_T_1088_data;
  assign T_1091 = T_1090[5:0];
  assign T_1095 = GEN_457 << tgtPages_T_1093_data;
  assign T_1096 = T_1095[5:0];
  assign T_1100 = GEN_457 << tgtPages_T_1098_data;
  assign T_1101 = T_1100[5:0];
  assign T_1105 = GEN_457 << tgtPages_T_1103_data;
  assign T_1106 = T_1105[5:0];
  assign T_1110 = GEN_457 << tgtPages_T_1108_data;
  assign T_1111 = T_1110[5:0];
  assign T_1115 = GEN_457 << tgtPages_T_1113_data;
  assign T_1116 = T_1115[5:0];
  assign T_1120 = GEN_457 << tgtPages_T_1118_data;
  assign T_1121 = T_1120[5:0];
  assign T_1125 = GEN_457 << tgtPages_T_1123_data;
  assign T_1126 = T_1125[5:0];
  assign T_1130 = GEN_457 << tgtPages_T_1128_data;
  assign T_1131 = T_1130[5:0];
  assign T_1135 = GEN_457 << tgtPages_T_1133_data;
  assign T_1136 = T_1135[5:0];
  assign T_1140 = GEN_457 << tgtPages_T_1138_data;
  assign T_1141 = T_1140[5:0];
  assign T_1145 = GEN_457 << tgtPages_T_1143_data;
  assign T_1146 = T_1145[5:0];
  assign T_1150 = GEN_457 << tgtPages_T_1148_data;
  assign T_1151 = T_1150[5:0];
  assign T_1155 = GEN_457 << tgtPages_T_1153_data;
  assign T_1156 = T_1155[5:0];
  assign T_1160 = GEN_457 << tgtPages_T_1158_data;
  assign T_1161 = T_1160[5:0];
  assign T_1165 = GEN_457 << tgtPages_T_1163_data;
  assign T_1166 = T_1165[5:0];
  assign T_1170 = GEN_457 << tgtPages_T_1168_data;
  assign T_1171 = T_1170[5:0];
  assign T_1175 = GEN_457 << tgtPages_T_1173_data;
  assign T_1176 = T_1175[5:0];
  assign T_1180 = GEN_457 << tgtPages_T_1178_data;
  assign T_1181 = T_1180[5:0];
  assign T_1185 = GEN_457 << tgtPages_T_1183_data;
  assign T_1186 = T_1185[5:0];
  assign T_1190 = GEN_457 << tgtPages_T_1188_data;
  assign T_1191 = T_1190[5:0];
  assign T_1195 = GEN_457 << tgtPages_T_1193_data;
  assign T_1196 = T_1195[5:0];
  assign brIdx_T_3612_addr = io_resp_bits_entry;
  assign brIdx_T_3612_en = 1'h1;
  `ifdef SYNTHESIS
  assign brIdx_T_3612_data = brIdx[brIdx_T_3612_addr];
  `else
  assign brIdx_T_3612_data = brIdx_T_3612_addr >= 6'h3e ? $random : brIdx[brIdx_T_3612_addr];
  `endif
  assign brIdx_T_2876_data = 1'h0;
  assign brIdx_T_2876_addr = T_2550;
  assign brIdx_T_2876_mask = r_btb_update_valid;
  assign brIdx_T_2876_en = r_btb_update_valid;
  assign GEN_4 = io_btb_update_valid ? io_btb_update_bits_prediction_valid : T_1216_prediction_valid;
  assign GEN_5 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_taken : T_1216_prediction_bits_taken;
  assign GEN_6 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_mask : T_1216_prediction_bits_mask;
  assign GEN_7 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bridx : T_1216_prediction_bits_bridx;
  assign GEN_8 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_target : T_1216_prediction_bits_target;
  assign GEN_9 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_entry : T_1216_prediction_bits_entry;
  assign GEN_10 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bht_history : T_1216_prediction_bits_bht_history;
  assign GEN_11 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bht_value : T_1216_prediction_bits_bht_value;
  assign GEN_12 = io_btb_update_valid ? io_btb_update_bits_pc : T_1216_pc;
  assign GEN_13 = io_btb_update_valid ? io_btb_update_bits_target : T_1216_target;
  assign GEN_14 = io_btb_update_valid ? io_btb_update_bits_taken : T_1216_taken;
  assign GEN_15 = io_btb_update_valid ? io_btb_update_bits_isJump : T_1216_isJump;
  assign GEN_16 = io_btb_update_valid ? io_btb_update_bits_isReturn : T_1216_isReturn;
  assign GEN_17 = io_btb_update_valid ? io_btb_update_bits_br_pc : T_1216_br_pc;
  assign r_btb_update_valid = T_1215;
  assign r_btb_update_bits_prediction_valid = T_1216_prediction_valid;
  assign r_btb_update_bits_prediction_bits_taken = T_1216_prediction_bits_taken;
  assign r_btb_update_bits_prediction_bits_mask = T_1216_prediction_bits_mask;
  assign r_btb_update_bits_prediction_bits_bridx = T_1216_prediction_bits_bridx;
  assign r_btb_update_bits_prediction_bits_target = T_1216_prediction_bits_target;
  assign r_btb_update_bits_prediction_bits_entry = T_1216_prediction_bits_entry;
  assign r_btb_update_bits_prediction_bits_bht_history = T_1216_prediction_bits_bht_history;
  assign r_btb_update_bits_prediction_bits_bht_value = T_1216_prediction_bits_bht_value;
  assign r_btb_update_bits_pc = T_1216_pc;
  assign r_btb_update_bits_target = T_1216_target;
  assign r_btb_update_bits_taken = T_1216_taken;
  assign r_btb_update_bits_isJump = T_1216_isJump;
  assign r_btb_update_bits_isReturn = T_1216_isReturn;
  assign r_btb_update_bits_br_pc = T_1216_br_pc;
  assign T_1398 = io_req_bits_addr[38:12];
  assign T_1401 = pages_T_1400_data == T_1398;
  assign T_1404 = pages_T_1403_data == T_1398;
  assign T_1407 = pages_T_1406_data == T_1398;
  assign T_1410 = pages_T_1409_data == T_1398;
  assign T_1413 = pages_T_1412_data == T_1398;
  assign T_1416 = pages_T_1415_data == T_1398;
  assign T_1422_0 = T_1401;
  assign T_1422_1 = T_1404;
  assign T_1422_2 = T_1407;
  assign T_1422_3 = T_1410;
  assign T_1422_4 = T_1413;
  assign T_1422_5 = T_1416;
  assign T_1424 = {T_1422_2,T_1422_1};
  assign T_1425 = {T_1424,T_1422_0};
  assign T_1426 = {T_1422_5,T_1422_4};
  assign T_1427 = {T_1426,T_1422_3};
  assign T_1428 = {T_1427,T_1425};
  assign pageHit = T_1428 & pageValid;
  assign T_1429 = io_req_bits_addr[11:0];
  assign T_1432 = idxs_T_1431_data == T_1429;
  assign T_1435 = idxs_T_1434_data == T_1429;
  assign T_1438 = idxs_T_1437_data == T_1429;
  assign T_1441 = idxs_T_1440_data == T_1429;
  assign T_1444 = idxs_T_1443_data == T_1429;
  assign T_1447 = idxs_T_1446_data == T_1429;
  assign T_1450 = idxs_T_1449_data == T_1429;
  assign T_1453 = idxs_T_1452_data == T_1429;
  assign T_1456 = idxs_T_1455_data == T_1429;
  assign T_1459 = idxs_T_1458_data == T_1429;
  assign T_1462 = idxs_T_1461_data == T_1429;
  assign T_1465 = idxs_T_1464_data == T_1429;
  assign T_1468 = idxs_T_1467_data == T_1429;
  assign T_1471 = idxs_T_1470_data == T_1429;
  assign T_1474 = idxs_T_1473_data == T_1429;
  assign T_1477 = idxs_T_1476_data == T_1429;
  assign T_1480 = idxs_T_1479_data == T_1429;
  assign T_1483 = idxs_T_1482_data == T_1429;
  assign T_1486 = idxs_T_1485_data == T_1429;
  assign T_1489 = idxs_T_1488_data == T_1429;
  assign T_1492 = idxs_T_1491_data == T_1429;
  assign T_1495 = idxs_T_1494_data == T_1429;
  assign T_1498 = idxs_T_1497_data == T_1429;
  assign T_1501 = idxs_T_1500_data == T_1429;
  assign T_1504 = idxs_T_1503_data == T_1429;
  assign T_1507 = idxs_T_1506_data == T_1429;
  assign T_1510 = idxs_T_1509_data == T_1429;
  assign T_1513 = idxs_T_1512_data == T_1429;
  assign T_1516 = idxs_T_1515_data == T_1429;
  assign T_1519 = idxs_T_1518_data == T_1429;
  assign T_1522 = idxs_T_1521_data == T_1429;
  assign T_1525 = idxs_T_1524_data == T_1429;
  assign T_1528 = idxs_T_1527_data == T_1429;
  assign T_1531 = idxs_T_1530_data == T_1429;
  assign T_1534 = idxs_T_1533_data == T_1429;
  assign T_1537 = idxs_T_1536_data == T_1429;
  assign T_1540 = idxs_T_1539_data == T_1429;
  assign T_1543 = idxs_T_1542_data == T_1429;
  assign T_1546 = idxs_T_1545_data == T_1429;
  assign T_1549 = idxs_T_1548_data == T_1429;
  assign T_1552 = idxs_T_1551_data == T_1429;
  assign T_1555 = idxs_T_1554_data == T_1429;
  assign T_1558 = idxs_T_1557_data == T_1429;
  assign T_1561 = idxs_T_1560_data == T_1429;
  assign T_1564 = idxs_T_1563_data == T_1429;
  assign T_1567 = idxs_T_1566_data == T_1429;
  assign T_1570 = idxs_T_1569_data == T_1429;
  assign T_1573 = idxs_T_1572_data == T_1429;
  assign T_1576 = idxs_T_1575_data == T_1429;
  assign T_1579 = idxs_T_1578_data == T_1429;
  assign T_1582 = idxs_T_1581_data == T_1429;
  assign T_1585 = idxs_T_1584_data == T_1429;
  assign T_1588 = idxs_T_1587_data == T_1429;
  assign T_1591 = idxs_T_1590_data == T_1429;
  assign T_1594 = idxs_T_1593_data == T_1429;
  assign T_1597 = idxs_T_1596_data == T_1429;
  assign T_1600 = idxs_T_1599_data == T_1429;
  assign T_1603 = idxs_T_1602_data == T_1429;
  assign T_1606 = idxs_T_1605_data == T_1429;
  assign T_1609 = idxs_T_1608_data == T_1429;
  assign T_1612 = idxs_T_1611_data == T_1429;
  assign T_1615 = idxs_T_1614_data == T_1429;
  assign T_1621_0 = T_1432;
  assign T_1621_1 = T_1435;
  assign T_1621_2 = T_1438;
  assign T_1621_3 = T_1441;
  assign T_1621_4 = T_1444;
  assign T_1621_5 = T_1447;
  assign T_1621_6 = T_1450;
  assign T_1621_7 = T_1453;
  assign T_1621_8 = T_1456;
  assign T_1621_9 = T_1459;
  assign T_1621_10 = T_1462;
  assign T_1621_11 = T_1465;
  assign T_1621_12 = T_1468;
  assign T_1621_13 = T_1471;
  assign T_1621_14 = T_1474;
  assign T_1621_15 = T_1477;
  assign T_1621_16 = T_1480;
  assign T_1621_17 = T_1483;
  assign T_1621_18 = T_1486;
  assign T_1621_19 = T_1489;
  assign T_1621_20 = T_1492;
  assign T_1621_21 = T_1495;
  assign T_1621_22 = T_1498;
  assign T_1621_23 = T_1501;
  assign T_1621_24 = T_1504;
  assign T_1621_25 = T_1507;
  assign T_1621_26 = T_1510;
  assign T_1621_27 = T_1513;
  assign T_1621_28 = T_1516;
  assign T_1621_29 = T_1519;
  assign T_1621_30 = T_1522;
  assign T_1621_31 = T_1525;
  assign T_1621_32 = T_1528;
  assign T_1621_33 = T_1531;
  assign T_1621_34 = T_1534;
  assign T_1621_35 = T_1537;
  assign T_1621_36 = T_1540;
  assign T_1621_37 = T_1543;
  assign T_1621_38 = T_1546;
  assign T_1621_39 = T_1549;
  assign T_1621_40 = T_1552;
  assign T_1621_41 = T_1555;
  assign T_1621_42 = T_1558;
  assign T_1621_43 = T_1561;
  assign T_1621_44 = T_1564;
  assign T_1621_45 = T_1567;
  assign T_1621_46 = T_1570;
  assign T_1621_47 = T_1573;
  assign T_1621_48 = T_1576;
  assign T_1621_49 = T_1579;
  assign T_1621_50 = T_1582;
  assign T_1621_51 = T_1585;
  assign T_1621_52 = T_1588;
  assign T_1621_53 = T_1591;
  assign T_1621_54 = T_1594;
  assign T_1621_55 = T_1597;
  assign T_1621_56 = T_1600;
  assign T_1621_57 = T_1603;
  assign T_1621_58 = T_1606;
  assign T_1621_59 = T_1609;
  assign T_1621_60 = T_1612;
  assign T_1621_61 = T_1615;
  assign T_1623 = {T_1621_2,T_1621_1};
  assign T_1624 = {T_1623,T_1621_0};
  assign T_1625 = {T_1621_4,T_1621_3};
  assign T_1626 = {T_1621_6,T_1621_5};
  assign T_1627 = {T_1626,T_1625};
  assign T_1628 = {T_1627,T_1624};
  assign T_1629 = {T_1621_8,T_1621_7};
  assign T_1630 = {T_1621_10,T_1621_9};
  assign T_1631 = {T_1630,T_1629};
  assign T_1632 = {T_1621_12,T_1621_11};
  assign T_1633 = {T_1621_14,T_1621_13};
  assign T_1634 = {T_1633,T_1632};
  assign T_1635 = {T_1634,T_1631};
  assign T_1636 = {T_1635,T_1628};
  assign T_1637 = {T_1621_16,T_1621_15};
  assign T_1638 = {T_1621_18,T_1621_17};
  assign T_1639 = {T_1638,T_1637};
  assign T_1640 = {T_1621_20,T_1621_19};
  assign T_1641 = {T_1621_22,T_1621_21};
  assign T_1642 = {T_1641,T_1640};
  assign T_1643 = {T_1642,T_1639};
  assign T_1644 = {T_1621_24,T_1621_23};
  assign T_1645 = {T_1621_26,T_1621_25};
  assign T_1646 = {T_1645,T_1644};
  assign T_1647 = {T_1621_28,T_1621_27};
  assign T_1648 = {T_1621_30,T_1621_29};
  assign T_1649 = {T_1648,T_1647};
  assign T_1650 = {T_1649,T_1646};
  assign T_1651 = {T_1650,T_1643};
  assign T_1652 = {T_1651,T_1636};
  assign T_1653 = {T_1621_33,T_1621_32};
  assign T_1654 = {T_1653,T_1621_31};
  assign T_1655 = {T_1621_35,T_1621_34};
  assign T_1656 = {T_1621_37,T_1621_36};
  assign T_1657 = {T_1656,T_1655};
  assign T_1658 = {T_1657,T_1654};
  assign T_1659 = {T_1621_39,T_1621_38};
  assign T_1660 = {T_1621_41,T_1621_40};
  assign T_1661 = {T_1660,T_1659};
  assign T_1662 = {T_1621_43,T_1621_42};
  assign T_1663 = {T_1621_45,T_1621_44};
  assign T_1664 = {T_1663,T_1662};
  assign T_1665 = {T_1664,T_1661};
  assign T_1666 = {T_1665,T_1658};
  assign T_1667 = {T_1621_47,T_1621_46};
  assign T_1668 = {T_1621_49,T_1621_48};
  assign T_1669 = {T_1668,T_1667};
  assign T_1670 = {T_1621_51,T_1621_50};
  assign T_1671 = {T_1621_53,T_1621_52};
  assign T_1672 = {T_1671,T_1670};
  assign T_1673 = {T_1672,T_1669};
  assign T_1674 = {T_1621_55,T_1621_54};
  assign T_1675 = {T_1621_57,T_1621_56};
  assign T_1676 = {T_1675,T_1674};
  assign T_1677 = {T_1621_59,T_1621_58};
  assign T_1678 = {T_1621_61,T_1621_60};
  assign T_1679 = {T_1678,T_1677};
  assign T_1680 = {T_1679,T_1676};
  assign T_1681 = {T_1680,T_1673};
  assign T_1682 = {T_1681,T_1666};
  assign T_1683 = {T_1682,T_1652};
  assign T_1684 = T_581 & pageHit;
  assign T_1685 = T_586 & pageHit;
  assign T_1686 = T_591 & pageHit;
  assign T_1687 = T_596 & pageHit;
  assign T_1688 = T_601 & pageHit;
  assign T_1689 = T_606 & pageHit;
  assign T_1690 = T_611 & pageHit;
  assign T_1691 = T_616 & pageHit;
  assign T_1692 = T_621 & pageHit;
  assign T_1693 = T_626 & pageHit;
  assign T_1694 = T_631 & pageHit;
  assign T_1695 = T_636 & pageHit;
  assign T_1696 = T_641 & pageHit;
  assign T_1697 = T_646 & pageHit;
  assign T_1698 = T_651 & pageHit;
  assign T_1699 = T_656 & pageHit;
  assign T_1700 = T_661 & pageHit;
  assign T_1701 = T_666 & pageHit;
  assign T_1702 = T_671 & pageHit;
  assign T_1703 = T_676 & pageHit;
  assign T_1704 = T_681 & pageHit;
  assign T_1705 = T_686 & pageHit;
  assign T_1706 = T_691 & pageHit;
  assign T_1707 = T_696 & pageHit;
  assign T_1708 = T_701 & pageHit;
  assign T_1709 = T_706 & pageHit;
  assign T_1710 = T_711 & pageHit;
  assign T_1711 = T_716 & pageHit;
  assign T_1712 = T_721 & pageHit;
  assign T_1713 = T_726 & pageHit;
  assign T_1714 = T_731 & pageHit;
  assign T_1715 = T_736 & pageHit;
  assign T_1716 = T_741 & pageHit;
  assign T_1717 = T_746 & pageHit;
  assign T_1718 = T_751 & pageHit;
  assign T_1719 = T_756 & pageHit;
  assign T_1720 = T_761 & pageHit;
  assign T_1721 = T_766 & pageHit;
  assign T_1722 = T_771 & pageHit;
  assign T_1723 = T_776 & pageHit;
  assign T_1724 = T_781 & pageHit;
  assign T_1725 = T_786 & pageHit;
  assign T_1726 = T_791 & pageHit;
  assign T_1727 = T_796 & pageHit;
  assign T_1728 = T_801 & pageHit;
  assign T_1729 = T_806 & pageHit;
  assign T_1730 = T_811 & pageHit;
  assign T_1731 = T_816 & pageHit;
  assign T_1732 = T_821 & pageHit;
  assign T_1733 = T_826 & pageHit;
  assign T_1734 = T_831 & pageHit;
  assign T_1735 = T_836 & pageHit;
  assign T_1736 = T_841 & pageHit;
  assign T_1737 = T_846 & pageHit;
  assign T_1738 = T_851 & pageHit;
  assign T_1739 = T_856 & pageHit;
  assign T_1740 = T_861 & pageHit;
  assign T_1741 = T_866 & pageHit;
  assign T_1742 = T_871 & pageHit;
  assign T_1743 = T_876 & pageHit;
  assign T_1744 = T_881 & pageHit;
  assign T_1745 = T_886 & pageHit;
  assign GEN_581 = {{5'd0}, 1'h0};
  assign T_1747 = T_1684 != GEN_581;
  assign T_1749 = T_1685 != GEN_581;
  assign T_1751 = T_1686 != GEN_581;
  assign T_1753 = T_1687 != GEN_581;
  assign T_1755 = T_1688 != GEN_581;
  assign T_1757 = T_1689 != GEN_581;
  assign T_1759 = T_1690 != GEN_581;
  assign T_1761 = T_1691 != GEN_581;
  assign T_1763 = T_1692 != GEN_581;
  assign T_1765 = T_1693 != GEN_581;
  assign T_1767 = T_1694 != GEN_581;
  assign T_1769 = T_1695 != GEN_581;
  assign T_1771 = T_1696 != GEN_581;
  assign T_1773 = T_1697 != GEN_581;
  assign T_1775 = T_1698 != GEN_581;
  assign T_1777 = T_1699 != GEN_581;
  assign T_1779 = T_1700 != GEN_581;
  assign T_1781 = T_1701 != GEN_581;
  assign T_1783 = T_1702 != GEN_581;
  assign T_1785 = T_1703 != GEN_581;
  assign T_1787 = T_1704 != GEN_581;
  assign T_1789 = T_1705 != GEN_581;
  assign T_1791 = T_1706 != GEN_581;
  assign T_1793 = T_1707 != GEN_581;
  assign T_1795 = T_1708 != GEN_581;
  assign T_1797 = T_1709 != GEN_581;
  assign T_1799 = T_1710 != GEN_581;
  assign T_1801 = T_1711 != GEN_581;
  assign T_1803 = T_1712 != GEN_581;
  assign T_1805 = T_1713 != GEN_581;
  assign T_1807 = T_1714 != GEN_581;
  assign T_1809 = T_1715 != GEN_581;
  assign T_1811 = T_1716 != GEN_581;
  assign T_1813 = T_1717 != GEN_581;
  assign T_1815 = T_1718 != GEN_581;
  assign T_1817 = T_1719 != GEN_581;
  assign T_1819 = T_1720 != GEN_581;
  assign T_1821 = T_1721 != GEN_581;
  assign T_1823 = T_1722 != GEN_581;
  assign T_1825 = T_1723 != GEN_581;
  assign T_1827 = T_1724 != GEN_581;
  assign T_1829 = T_1725 != GEN_581;
  assign T_1831 = T_1726 != GEN_581;
  assign T_1833 = T_1727 != GEN_581;
  assign T_1835 = T_1728 != GEN_581;
  assign T_1837 = T_1729 != GEN_581;
  assign T_1839 = T_1730 != GEN_581;
  assign T_1841 = T_1731 != GEN_581;
  assign T_1843 = T_1732 != GEN_581;
  assign T_1845 = T_1733 != GEN_581;
  assign T_1847 = T_1734 != GEN_581;
  assign T_1849 = T_1735 != GEN_581;
  assign T_1851 = T_1736 != GEN_581;
  assign T_1853 = T_1737 != GEN_581;
  assign T_1855 = T_1738 != GEN_581;
  assign T_1857 = T_1739 != GEN_581;
  assign T_1859 = T_1740 != GEN_581;
  assign T_1861 = T_1741 != GEN_581;
  assign T_1863 = T_1742 != GEN_581;
  assign T_1865 = T_1743 != GEN_581;
  assign T_1867 = T_1744 != GEN_581;
  assign T_1869 = T_1745 != GEN_581;
  assign T_1875_0 = T_1747;
  assign T_1875_1 = T_1749;
  assign T_1875_2 = T_1751;
  assign T_1875_3 = T_1753;
  assign T_1875_4 = T_1755;
  assign T_1875_5 = T_1757;
  assign T_1875_6 = T_1759;
  assign T_1875_7 = T_1761;
  assign T_1875_8 = T_1763;
  assign T_1875_9 = T_1765;
  assign T_1875_10 = T_1767;
  assign T_1875_11 = T_1769;
  assign T_1875_12 = T_1771;
  assign T_1875_13 = T_1773;
  assign T_1875_14 = T_1775;
  assign T_1875_15 = T_1777;
  assign T_1875_16 = T_1779;
  assign T_1875_17 = T_1781;
  assign T_1875_18 = T_1783;
  assign T_1875_19 = T_1785;
  assign T_1875_20 = T_1787;
  assign T_1875_21 = T_1789;
  assign T_1875_22 = T_1791;
  assign T_1875_23 = T_1793;
  assign T_1875_24 = T_1795;
  assign T_1875_25 = T_1797;
  assign T_1875_26 = T_1799;
  assign T_1875_27 = T_1801;
  assign T_1875_28 = T_1803;
  assign T_1875_29 = T_1805;
  assign T_1875_30 = T_1807;
  assign T_1875_31 = T_1809;
  assign T_1875_32 = T_1811;
  assign T_1875_33 = T_1813;
  assign T_1875_34 = T_1815;
  assign T_1875_35 = T_1817;
  assign T_1875_36 = T_1819;
  assign T_1875_37 = T_1821;
  assign T_1875_38 = T_1823;
  assign T_1875_39 = T_1825;
  assign T_1875_40 = T_1827;
  assign T_1875_41 = T_1829;
  assign T_1875_42 = T_1831;
  assign T_1875_43 = T_1833;
  assign T_1875_44 = T_1835;
  assign T_1875_45 = T_1837;
  assign T_1875_46 = T_1839;
  assign T_1875_47 = T_1841;
  assign T_1875_48 = T_1843;
  assign T_1875_49 = T_1845;
  assign T_1875_50 = T_1847;
  assign T_1875_51 = T_1849;
  assign T_1875_52 = T_1851;
  assign T_1875_53 = T_1853;
  assign T_1875_54 = T_1855;
  assign T_1875_55 = T_1857;
  assign T_1875_56 = T_1859;
  assign T_1875_57 = T_1861;
  assign T_1875_58 = T_1863;
  assign T_1875_59 = T_1865;
  assign T_1875_60 = T_1867;
  assign T_1875_61 = T_1869;
  assign T_1877 = {T_1875_2,T_1875_1};
  assign T_1878 = {T_1877,T_1875_0};
  assign T_1879 = {T_1875_4,T_1875_3};
  assign T_1880 = {T_1875_6,T_1875_5};
  assign T_1881 = {T_1880,T_1879};
  assign T_1882 = {T_1881,T_1878};
  assign T_1883 = {T_1875_8,T_1875_7};
  assign T_1884 = {T_1875_10,T_1875_9};
  assign T_1885 = {T_1884,T_1883};
  assign T_1886 = {T_1875_12,T_1875_11};
  assign T_1887 = {T_1875_14,T_1875_13};
  assign T_1888 = {T_1887,T_1886};
  assign T_1889 = {T_1888,T_1885};
  assign T_1890 = {T_1889,T_1882};
  assign T_1891 = {T_1875_16,T_1875_15};
  assign T_1892 = {T_1875_18,T_1875_17};
  assign T_1893 = {T_1892,T_1891};
  assign T_1894 = {T_1875_20,T_1875_19};
  assign T_1895 = {T_1875_22,T_1875_21};
  assign T_1896 = {T_1895,T_1894};
  assign T_1897 = {T_1896,T_1893};
  assign T_1898 = {T_1875_24,T_1875_23};
  assign T_1899 = {T_1875_26,T_1875_25};
  assign T_1900 = {T_1899,T_1898};
  assign T_1901 = {T_1875_28,T_1875_27};
  assign T_1902 = {T_1875_30,T_1875_29};
  assign T_1903 = {T_1902,T_1901};
  assign T_1904 = {T_1903,T_1900};
  assign T_1905 = {T_1904,T_1897};
  assign T_1906 = {T_1905,T_1890};
  assign T_1907 = {T_1875_33,T_1875_32};
  assign T_1908 = {T_1907,T_1875_31};
  assign T_1909 = {T_1875_35,T_1875_34};
  assign T_1910 = {T_1875_37,T_1875_36};
  assign T_1911 = {T_1910,T_1909};
  assign T_1912 = {T_1911,T_1908};
  assign T_1913 = {T_1875_39,T_1875_38};
  assign T_1914 = {T_1875_41,T_1875_40};
  assign T_1915 = {T_1914,T_1913};
  assign T_1916 = {T_1875_43,T_1875_42};
  assign T_1917 = {T_1875_45,T_1875_44};
  assign T_1918 = {T_1917,T_1916};
  assign T_1919 = {T_1918,T_1915};
  assign T_1920 = {T_1919,T_1912};
  assign T_1921 = {T_1875_47,T_1875_46};
  assign T_1922 = {T_1875_49,T_1875_48};
  assign T_1923 = {T_1922,T_1921};
  assign T_1924 = {T_1875_51,T_1875_50};
  assign T_1925 = {T_1875_53,T_1875_52};
  assign T_1926 = {T_1925,T_1924};
  assign T_1927 = {T_1926,T_1923};
  assign T_1928 = {T_1875_55,T_1875_54};
  assign T_1929 = {T_1875_57,T_1875_56};
  assign T_1930 = {T_1929,T_1928};
  assign T_1931 = {T_1875_59,T_1875_58};
  assign T_1932 = {T_1875_61,T_1875_60};
  assign T_1933 = {T_1932,T_1931};
  assign T_1934 = {T_1933,T_1930};
  assign T_1935 = {T_1934,T_1927};
  assign T_1936 = {T_1935,T_1920};
  assign T_1937 = {T_1936,T_1906};
  assign T_1938 = idxValid & T_1683;
  assign hits = T_1938 & T_1937;
  assign T_1939 = r_btb_update_bits_pc[38:12];
  assign T_1942 = pages_T_1941_data == T_1939;
  assign T_1945 = pages_T_1944_data == T_1939;
  assign T_1948 = pages_T_1947_data == T_1939;
  assign T_1951 = pages_T_1950_data == T_1939;
  assign T_1954 = pages_T_1953_data == T_1939;
  assign T_1957 = pages_T_1956_data == T_1939;
  assign T_1963_0 = T_1942;
  assign T_1963_1 = T_1945;
  assign T_1963_2 = T_1948;
  assign T_1963_3 = T_1951;
  assign T_1963_4 = T_1954;
  assign T_1963_5 = T_1957;
  assign T_1965 = {T_1963_2,T_1963_1};
  assign T_1966 = {T_1965,T_1963_0};
  assign T_1967 = {T_1963_5,T_1963_4};
  assign T_1968 = {T_1967,T_1963_3};
  assign T_1969 = {T_1968,T_1966};
  assign updatePageHit = T_1969 & pageValid;
  assign T_1970 = r_btb_update_bits_pc[11:0];
  assign T_1973 = idxs_T_1972_data == T_1970;
  assign T_1976 = idxs_T_1975_data == T_1970;
  assign T_1979 = idxs_T_1978_data == T_1970;
  assign T_1982 = idxs_T_1981_data == T_1970;
  assign T_1985 = idxs_T_1984_data == T_1970;
  assign T_1988 = idxs_T_1987_data == T_1970;
  assign T_1991 = idxs_T_1990_data == T_1970;
  assign T_1994 = idxs_T_1993_data == T_1970;
  assign T_1997 = idxs_T_1996_data == T_1970;
  assign T_2000 = idxs_T_1999_data == T_1970;
  assign T_2003 = idxs_T_2002_data == T_1970;
  assign T_2006 = idxs_T_2005_data == T_1970;
  assign T_2009 = idxs_T_2008_data == T_1970;
  assign T_2012 = idxs_T_2011_data == T_1970;
  assign T_2015 = idxs_T_2014_data == T_1970;
  assign T_2018 = idxs_T_2017_data == T_1970;
  assign T_2021 = idxs_T_2020_data == T_1970;
  assign T_2024 = idxs_T_2023_data == T_1970;
  assign T_2027 = idxs_T_2026_data == T_1970;
  assign T_2030 = idxs_T_2029_data == T_1970;
  assign T_2033 = idxs_T_2032_data == T_1970;
  assign T_2036 = idxs_T_2035_data == T_1970;
  assign T_2039 = idxs_T_2038_data == T_1970;
  assign T_2042 = idxs_T_2041_data == T_1970;
  assign T_2045 = idxs_T_2044_data == T_1970;
  assign T_2048 = idxs_T_2047_data == T_1970;
  assign T_2051 = idxs_T_2050_data == T_1970;
  assign T_2054 = idxs_T_2053_data == T_1970;
  assign T_2057 = idxs_T_2056_data == T_1970;
  assign T_2060 = idxs_T_2059_data == T_1970;
  assign T_2063 = idxs_T_2062_data == T_1970;
  assign T_2066 = idxs_T_2065_data == T_1970;
  assign T_2069 = idxs_T_2068_data == T_1970;
  assign T_2072 = idxs_T_2071_data == T_1970;
  assign T_2075 = idxs_T_2074_data == T_1970;
  assign T_2078 = idxs_T_2077_data == T_1970;
  assign T_2081 = idxs_T_2080_data == T_1970;
  assign T_2084 = idxs_T_2083_data == T_1970;
  assign T_2087 = idxs_T_2086_data == T_1970;
  assign T_2090 = idxs_T_2089_data == T_1970;
  assign T_2093 = idxs_T_2092_data == T_1970;
  assign T_2096 = idxs_T_2095_data == T_1970;
  assign T_2099 = idxs_T_2098_data == T_1970;
  assign T_2102 = idxs_T_2101_data == T_1970;
  assign T_2105 = idxs_T_2104_data == T_1970;
  assign T_2108 = idxs_T_2107_data == T_1970;
  assign T_2111 = idxs_T_2110_data == T_1970;
  assign T_2114 = idxs_T_2113_data == T_1970;
  assign T_2117 = idxs_T_2116_data == T_1970;
  assign T_2120 = idxs_T_2119_data == T_1970;
  assign T_2123 = idxs_T_2122_data == T_1970;
  assign T_2126 = idxs_T_2125_data == T_1970;
  assign T_2129 = idxs_T_2128_data == T_1970;
  assign T_2132 = idxs_T_2131_data == T_1970;
  assign T_2135 = idxs_T_2134_data == T_1970;
  assign T_2138 = idxs_T_2137_data == T_1970;
  assign T_2141 = idxs_T_2140_data == T_1970;
  assign T_2144 = idxs_T_2143_data == T_1970;
  assign T_2147 = idxs_T_2146_data == T_1970;
  assign T_2150 = idxs_T_2149_data == T_1970;
  assign T_2153 = idxs_T_2152_data == T_1970;
  assign T_2156 = idxs_T_2155_data == T_1970;
  assign T_2162_0 = T_1973;
  assign T_2162_1 = T_1976;
  assign T_2162_2 = T_1979;
  assign T_2162_3 = T_1982;
  assign T_2162_4 = T_1985;
  assign T_2162_5 = T_1988;
  assign T_2162_6 = T_1991;
  assign T_2162_7 = T_1994;
  assign T_2162_8 = T_1997;
  assign T_2162_9 = T_2000;
  assign T_2162_10 = T_2003;
  assign T_2162_11 = T_2006;
  assign T_2162_12 = T_2009;
  assign T_2162_13 = T_2012;
  assign T_2162_14 = T_2015;
  assign T_2162_15 = T_2018;
  assign T_2162_16 = T_2021;
  assign T_2162_17 = T_2024;
  assign T_2162_18 = T_2027;
  assign T_2162_19 = T_2030;
  assign T_2162_20 = T_2033;
  assign T_2162_21 = T_2036;
  assign T_2162_22 = T_2039;
  assign T_2162_23 = T_2042;
  assign T_2162_24 = T_2045;
  assign T_2162_25 = T_2048;
  assign T_2162_26 = T_2051;
  assign T_2162_27 = T_2054;
  assign T_2162_28 = T_2057;
  assign T_2162_29 = T_2060;
  assign T_2162_30 = T_2063;
  assign T_2162_31 = T_2066;
  assign T_2162_32 = T_2069;
  assign T_2162_33 = T_2072;
  assign T_2162_34 = T_2075;
  assign T_2162_35 = T_2078;
  assign T_2162_36 = T_2081;
  assign T_2162_37 = T_2084;
  assign T_2162_38 = T_2087;
  assign T_2162_39 = T_2090;
  assign T_2162_40 = T_2093;
  assign T_2162_41 = T_2096;
  assign T_2162_42 = T_2099;
  assign T_2162_43 = T_2102;
  assign T_2162_44 = T_2105;
  assign T_2162_45 = T_2108;
  assign T_2162_46 = T_2111;
  assign T_2162_47 = T_2114;
  assign T_2162_48 = T_2117;
  assign T_2162_49 = T_2120;
  assign T_2162_50 = T_2123;
  assign T_2162_51 = T_2126;
  assign T_2162_52 = T_2129;
  assign T_2162_53 = T_2132;
  assign T_2162_54 = T_2135;
  assign T_2162_55 = T_2138;
  assign T_2162_56 = T_2141;
  assign T_2162_57 = T_2144;
  assign T_2162_58 = T_2147;
  assign T_2162_59 = T_2150;
  assign T_2162_60 = T_2153;
  assign T_2162_61 = T_2156;
  assign T_2225 = T_581 & updatePageHit;
  assign T_2226 = T_586 & updatePageHit;
  assign T_2227 = T_591 & updatePageHit;
  assign T_2228 = T_596 & updatePageHit;
  assign T_2229 = T_601 & updatePageHit;
  assign T_2230 = T_606 & updatePageHit;
  assign T_2231 = T_611 & updatePageHit;
  assign T_2232 = T_616 & updatePageHit;
  assign T_2233 = T_621 & updatePageHit;
  assign T_2234 = T_626 & updatePageHit;
  assign T_2235 = T_631 & updatePageHit;
  assign T_2236 = T_636 & updatePageHit;
  assign T_2237 = T_641 & updatePageHit;
  assign T_2238 = T_646 & updatePageHit;
  assign T_2239 = T_651 & updatePageHit;
  assign T_2240 = T_656 & updatePageHit;
  assign T_2241 = T_661 & updatePageHit;
  assign T_2242 = T_666 & updatePageHit;
  assign T_2243 = T_671 & updatePageHit;
  assign T_2244 = T_676 & updatePageHit;
  assign T_2245 = T_681 & updatePageHit;
  assign T_2246 = T_686 & updatePageHit;
  assign T_2247 = T_691 & updatePageHit;
  assign T_2248 = T_696 & updatePageHit;
  assign T_2249 = T_701 & updatePageHit;
  assign T_2250 = T_706 & updatePageHit;
  assign T_2251 = T_711 & updatePageHit;
  assign T_2252 = T_716 & updatePageHit;
  assign T_2253 = T_721 & updatePageHit;
  assign T_2254 = T_726 & updatePageHit;
  assign T_2255 = T_731 & updatePageHit;
  assign T_2256 = T_736 & updatePageHit;
  assign T_2257 = T_741 & updatePageHit;
  assign T_2258 = T_746 & updatePageHit;
  assign T_2259 = T_751 & updatePageHit;
  assign T_2260 = T_756 & updatePageHit;
  assign T_2261 = T_761 & updatePageHit;
  assign T_2262 = T_766 & updatePageHit;
  assign T_2263 = T_771 & updatePageHit;
  assign T_2264 = T_776 & updatePageHit;
  assign T_2265 = T_781 & updatePageHit;
  assign T_2266 = T_786 & updatePageHit;
  assign T_2267 = T_791 & updatePageHit;
  assign T_2268 = T_796 & updatePageHit;
  assign T_2269 = T_801 & updatePageHit;
  assign T_2270 = T_806 & updatePageHit;
  assign T_2271 = T_811 & updatePageHit;
  assign T_2272 = T_816 & updatePageHit;
  assign T_2273 = T_821 & updatePageHit;
  assign T_2274 = T_826 & updatePageHit;
  assign T_2275 = T_831 & updatePageHit;
  assign T_2276 = T_836 & updatePageHit;
  assign T_2277 = T_841 & updatePageHit;
  assign T_2278 = T_846 & updatePageHit;
  assign T_2279 = T_851 & updatePageHit;
  assign T_2280 = T_856 & updatePageHit;
  assign T_2281 = T_861 & updatePageHit;
  assign T_2282 = T_866 & updatePageHit;
  assign T_2283 = T_871 & updatePageHit;
  assign T_2284 = T_876 & updatePageHit;
  assign T_2285 = T_881 & updatePageHit;
  assign T_2286 = T_886 & updatePageHit;
  assign T_2288 = T_2225 != GEN_581;
  assign T_2290 = T_2226 != GEN_581;
  assign T_2292 = T_2227 != GEN_581;
  assign T_2294 = T_2228 != GEN_581;
  assign T_2296 = T_2229 != GEN_581;
  assign T_2298 = T_2230 != GEN_581;
  assign T_2300 = T_2231 != GEN_581;
  assign T_2302 = T_2232 != GEN_581;
  assign T_2304 = T_2233 != GEN_581;
  assign T_2306 = T_2234 != GEN_581;
  assign T_2308 = T_2235 != GEN_581;
  assign T_2310 = T_2236 != GEN_581;
  assign T_2312 = T_2237 != GEN_581;
  assign T_2314 = T_2238 != GEN_581;
  assign T_2316 = T_2239 != GEN_581;
  assign T_2318 = T_2240 != GEN_581;
  assign T_2320 = T_2241 != GEN_581;
  assign T_2322 = T_2242 != GEN_581;
  assign T_2324 = T_2243 != GEN_581;
  assign T_2326 = T_2244 != GEN_581;
  assign T_2328 = T_2245 != GEN_581;
  assign T_2330 = T_2246 != GEN_581;
  assign T_2332 = T_2247 != GEN_581;
  assign T_2334 = T_2248 != GEN_581;
  assign T_2336 = T_2249 != GEN_581;
  assign T_2338 = T_2250 != GEN_581;
  assign T_2340 = T_2251 != GEN_581;
  assign T_2342 = T_2252 != GEN_581;
  assign T_2344 = T_2253 != GEN_581;
  assign T_2346 = T_2254 != GEN_581;
  assign T_2348 = T_2255 != GEN_581;
  assign T_2350 = T_2256 != GEN_581;
  assign T_2352 = T_2257 != GEN_581;
  assign T_2354 = T_2258 != GEN_581;
  assign T_2356 = T_2259 != GEN_581;
  assign T_2358 = T_2260 != GEN_581;
  assign T_2360 = T_2261 != GEN_581;
  assign T_2362 = T_2262 != GEN_581;
  assign T_2364 = T_2263 != GEN_581;
  assign T_2366 = T_2264 != GEN_581;
  assign T_2368 = T_2265 != GEN_581;
  assign T_2370 = T_2266 != GEN_581;
  assign T_2372 = T_2267 != GEN_581;
  assign T_2374 = T_2268 != GEN_581;
  assign T_2376 = T_2269 != GEN_581;
  assign T_2378 = T_2270 != GEN_581;
  assign T_2380 = T_2271 != GEN_581;
  assign T_2382 = T_2272 != GEN_581;
  assign T_2384 = T_2273 != GEN_581;
  assign T_2386 = T_2274 != GEN_581;
  assign T_2388 = T_2275 != GEN_581;
  assign T_2390 = T_2276 != GEN_581;
  assign T_2392 = T_2277 != GEN_581;
  assign T_2394 = T_2278 != GEN_581;
  assign T_2396 = T_2279 != GEN_581;
  assign T_2398 = T_2280 != GEN_581;
  assign T_2400 = T_2281 != GEN_581;
  assign T_2402 = T_2282 != GEN_581;
  assign T_2404 = T_2283 != GEN_581;
  assign T_2406 = T_2284 != GEN_581;
  assign T_2408 = T_2285 != GEN_581;
  assign T_2410 = T_2286 != GEN_581;
  assign T_2416_0 = T_2288;
  assign T_2416_1 = T_2290;
  assign T_2416_2 = T_2292;
  assign T_2416_3 = T_2294;
  assign T_2416_4 = T_2296;
  assign T_2416_5 = T_2298;
  assign T_2416_6 = T_2300;
  assign T_2416_7 = T_2302;
  assign T_2416_8 = T_2304;
  assign T_2416_9 = T_2306;
  assign T_2416_10 = T_2308;
  assign T_2416_11 = T_2310;
  assign T_2416_12 = T_2312;
  assign T_2416_13 = T_2314;
  assign T_2416_14 = T_2316;
  assign T_2416_15 = T_2318;
  assign T_2416_16 = T_2320;
  assign T_2416_17 = T_2322;
  assign T_2416_18 = T_2324;
  assign T_2416_19 = T_2326;
  assign T_2416_20 = T_2328;
  assign T_2416_21 = T_2330;
  assign T_2416_22 = T_2332;
  assign T_2416_23 = T_2334;
  assign T_2416_24 = T_2336;
  assign T_2416_25 = T_2338;
  assign T_2416_26 = T_2340;
  assign T_2416_27 = T_2342;
  assign T_2416_28 = T_2344;
  assign T_2416_29 = T_2346;
  assign T_2416_30 = T_2348;
  assign T_2416_31 = T_2350;
  assign T_2416_32 = T_2352;
  assign T_2416_33 = T_2354;
  assign T_2416_34 = T_2356;
  assign T_2416_35 = T_2358;
  assign T_2416_36 = T_2360;
  assign T_2416_37 = T_2362;
  assign T_2416_38 = T_2364;
  assign T_2416_39 = T_2366;
  assign T_2416_40 = T_2368;
  assign T_2416_41 = T_2370;
  assign T_2416_42 = T_2372;
  assign T_2416_43 = T_2374;
  assign T_2416_44 = T_2376;
  assign T_2416_45 = T_2378;
  assign T_2416_46 = T_2380;
  assign T_2416_47 = T_2382;
  assign T_2416_48 = T_2384;
  assign T_2416_49 = T_2386;
  assign T_2416_50 = T_2388;
  assign T_2416_51 = T_2390;
  assign T_2416_52 = T_2392;
  assign T_2416_53 = T_2394;
  assign T_2416_54 = T_2396;
  assign T_2416_55 = T_2398;
  assign T_2416_56 = T_2400;
  assign T_2416_57 = T_2402;
  assign T_2416_58 = T_2404;
  assign T_2416_59 = T_2406;
  assign T_2416_60 = T_2408;
  assign T_2416_61 = T_2410;
  assign T_2481 = r_btb_update_bits_prediction_valid == 1'h0;
  assign T_2482 = r_btb_update_valid & T_2481;
  assign T_2485 = nextRepl == 6'h3d;
  assign GEN_705 = {{5'd0}, 1'h1};
  assign T_2487 = nextRepl + GEN_705;
  assign T_2488 = T_2487[5:0];
  assign GEN_18 = T_2485 ? {{5'd0}, 1'h0} : T_2488;
  assign GEN_19 = T_2482 ? GEN_18 : nextRepl;
  assign useUpdatePageHit = updatePageHit != GEN_581;
  assign doIdxPageRepl = useUpdatePageHit == 1'h0;
  assign idxPageRepl = T_2545[5:0];
  assign idxPageUpdateOH = useUpdatePageHit ? updatePageHit : idxPageRepl;
  assign T_2494 = idxPageUpdateOH[5:4];
  assign T_2495 = idxPageUpdateOH[3:0];
  assign GEN_707 = {{1'd0}, 1'h0};
  assign T_2497 = T_2494 != GEN_707;
  assign GEN_708 = {{2'd0}, T_2494};
  assign T_2498 = GEN_708 | T_2495;
  assign T_2499 = T_2498[3:2];
  assign T_2500 = T_2498[1:0];
  assign T_2502 = T_2499 != GEN_707;
  assign T_2503 = T_2499 | T_2500;
  assign T_2504 = T_2503[1];
  assign T_2505 = {T_2502,T_2504};
  assign idxPageUpdate = {T_2497,T_2505};
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : {{5'd0}, 1'h0};
  assign samePage = T_1939 == T_1398;
  assign T_2509 = ~ idxPageReplEn;
  assign T_2510 = pageHit & T_2509;
  assign usePageHit = T_2510 != GEN_581;
  assign T_2513 = samePage == 1'h0;
  assign T_2515 = usePageHit == 1'h0;
  assign doTgtPageRepl = T_2513 & T_2515;
  assign T_2516 = idxPageUpdateOH[4:0];
  assign GEN_711 = {{1'd0}, T_2516};
  assign T_2517 = GEN_711 << 1;
  assign T_2518 = idxPageUpdateOH[5];
  assign GEN_712 = {{5'd0}, T_2518};
  assign T_2519 = T_2517 | GEN_712;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T_2519;
  assign T_2520 = usePageHit ? pageHit : tgtPageRepl;
  assign T_2521 = T_2520[5:4];
  assign T_2522 = T_2520[3:0];
  assign T_2524 = T_2521 != GEN_707;
  assign GEN_714 = {{2'd0}, T_2521};
  assign T_2525 = GEN_714 | T_2522;
  assign T_2526 = T_2525[3:2];
  assign T_2527 = T_2525[1:0];
  assign T_2529 = T_2526 != GEN_707;
  assign T_2530 = T_2526 | T_2527;
  assign T_2531 = T_2530[1];
  assign T_2532 = {T_2529,T_2531};
  assign tgtPageUpdate = {T_2524,T_2532};
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : {{5'd0}, 1'h0};
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign T_2534 = r_btb_update_valid & doPageRepl;
  assign T_2538 = T_2536 == 3'h5;
  assign GEN_716 = {{2'd0}, 1'h1};
  assign T_2540 = T_2536 + GEN_716;
  assign T_2541 = T_2540[2:0];
  assign GEN_20 = T_2538 ? {{2'd0}, 1'h0} : T_2541;
  assign GEN_21 = T_2534 ? GEN_20 : T_2536;
  assign T_2545 = GEN_457 << T_2536;
  assign T_2546 = io_req_bits_addr == r_btb_update_bits_target;
  assign T_2547 = T_2546 | reset;
  assign T_2549 = T_2547 == 1'h0;
  assign T_2550 = r_btb_update_bits_prediction_valid ? r_btb_update_bits_prediction_bits_entry : nextRepl;
  assign T_2551 = T_581 | T_891;
  assign T_2552 = pageReplEn & T_2551;
  assign T_2554 = T_2552 != GEN_581;
  assign T_2555 = T_586 | T_896;
  assign T_2556 = pageReplEn & T_2555;
  assign T_2558 = T_2556 != GEN_581;
  assign T_2559 = T_591 | T_901;
  assign T_2560 = pageReplEn & T_2559;
  assign T_2562 = T_2560 != GEN_581;
  assign T_2563 = T_596 | T_906;
  assign T_2564 = pageReplEn & T_2563;
  assign T_2566 = T_2564 != GEN_581;
  assign T_2567 = T_601 | T_911;
  assign T_2568 = pageReplEn & T_2567;
  assign T_2570 = T_2568 != GEN_581;
  assign T_2571 = T_606 | T_916;
  assign T_2572 = pageReplEn & T_2571;
  assign T_2574 = T_2572 != GEN_581;
  assign T_2575 = T_611 | T_921;
  assign T_2576 = pageReplEn & T_2575;
  assign T_2578 = T_2576 != GEN_581;
  assign T_2579 = T_616 | T_926;
  assign T_2580 = pageReplEn & T_2579;
  assign T_2582 = T_2580 != GEN_581;
  assign T_2583 = T_621 | T_931;
  assign T_2584 = pageReplEn & T_2583;
  assign T_2586 = T_2584 != GEN_581;
  assign T_2587 = T_626 | T_936;
  assign T_2588 = pageReplEn & T_2587;
  assign T_2590 = T_2588 != GEN_581;
  assign T_2591 = T_631 | T_941;
  assign T_2592 = pageReplEn & T_2591;
  assign T_2594 = T_2592 != GEN_581;
  assign T_2595 = T_636 | T_946;
  assign T_2596 = pageReplEn & T_2595;
  assign T_2598 = T_2596 != GEN_581;
  assign T_2599 = T_641 | T_951;
  assign T_2600 = pageReplEn & T_2599;
  assign T_2602 = T_2600 != GEN_581;
  assign T_2603 = T_646 | T_956;
  assign T_2604 = pageReplEn & T_2603;
  assign T_2606 = T_2604 != GEN_581;
  assign T_2607 = T_651 | T_961;
  assign T_2608 = pageReplEn & T_2607;
  assign T_2610 = T_2608 != GEN_581;
  assign T_2611 = T_656 | T_966;
  assign T_2612 = pageReplEn & T_2611;
  assign T_2614 = T_2612 != GEN_581;
  assign T_2615 = T_661 | T_971;
  assign T_2616 = pageReplEn & T_2615;
  assign T_2618 = T_2616 != GEN_581;
  assign T_2619 = T_666 | T_976;
  assign T_2620 = pageReplEn & T_2619;
  assign T_2622 = T_2620 != GEN_581;
  assign T_2623 = T_671 | T_981;
  assign T_2624 = pageReplEn & T_2623;
  assign T_2626 = T_2624 != GEN_581;
  assign T_2627 = T_676 | T_986;
  assign T_2628 = pageReplEn & T_2627;
  assign T_2630 = T_2628 != GEN_581;
  assign T_2631 = T_681 | T_991;
  assign T_2632 = pageReplEn & T_2631;
  assign T_2634 = T_2632 != GEN_581;
  assign T_2635 = T_686 | T_996;
  assign T_2636 = pageReplEn & T_2635;
  assign T_2638 = T_2636 != GEN_581;
  assign T_2639 = T_691 | T_1001;
  assign T_2640 = pageReplEn & T_2639;
  assign T_2642 = T_2640 != GEN_581;
  assign T_2643 = T_696 | T_1006;
  assign T_2644 = pageReplEn & T_2643;
  assign T_2646 = T_2644 != GEN_581;
  assign T_2647 = T_701 | T_1011;
  assign T_2648 = pageReplEn & T_2647;
  assign T_2650 = T_2648 != GEN_581;
  assign T_2651 = T_706 | T_1016;
  assign T_2652 = pageReplEn & T_2651;
  assign T_2654 = T_2652 != GEN_581;
  assign T_2655 = T_711 | T_1021;
  assign T_2656 = pageReplEn & T_2655;
  assign T_2658 = T_2656 != GEN_581;
  assign T_2659 = T_716 | T_1026;
  assign T_2660 = pageReplEn & T_2659;
  assign T_2662 = T_2660 != GEN_581;
  assign T_2663 = T_721 | T_1031;
  assign T_2664 = pageReplEn & T_2663;
  assign T_2666 = T_2664 != GEN_581;
  assign T_2667 = T_726 | T_1036;
  assign T_2668 = pageReplEn & T_2667;
  assign T_2670 = T_2668 != GEN_581;
  assign T_2671 = T_731 | T_1041;
  assign T_2672 = pageReplEn & T_2671;
  assign T_2674 = T_2672 != GEN_581;
  assign T_2675 = T_736 | T_1046;
  assign T_2676 = pageReplEn & T_2675;
  assign T_2678 = T_2676 != GEN_581;
  assign T_2679 = T_741 | T_1051;
  assign T_2680 = pageReplEn & T_2679;
  assign T_2682 = T_2680 != GEN_581;
  assign T_2683 = T_746 | T_1056;
  assign T_2684 = pageReplEn & T_2683;
  assign T_2686 = T_2684 != GEN_581;
  assign T_2687 = T_751 | T_1061;
  assign T_2688 = pageReplEn & T_2687;
  assign T_2690 = T_2688 != GEN_581;
  assign T_2691 = T_756 | T_1066;
  assign T_2692 = pageReplEn & T_2691;
  assign T_2694 = T_2692 != GEN_581;
  assign T_2695 = T_761 | T_1071;
  assign T_2696 = pageReplEn & T_2695;
  assign T_2698 = T_2696 != GEN_581;
  assign T_2699 = T_766 | T_1076;
  assign T_2700 = pageReplEn & T_2699;
  assign T_2702 = T_2700 != GEN_581;
  assign T_2703 = T_771 | T_1081;
  assign T_2704 = pageReplEn & T_2703;
  assign T_2706 = T_2704 != GEN_581;
  assign T_2707 = T_776 | T_1086;
  assign T_2708 = pageReplEn & T_2707;
  assign T_2710 = T_2708 != GEN_581;
  assign T_2711 = T_781 | T_1091;
  assign T_2712 = pageReplEn & T_2711;
  assign T_2714 = T_2712 != GEN_581;
  assign T_2715 = T_786 | T_1096;
  assign T_2716 = pageReplEn & T_2715;
  assign T_2718 = T_2716 != GEN_581;
  assign T_2719 = T_791 | T_1101;
  assign T_2720 = pageReplEn & T_2719;
  assign T_2722 = T_2720 != GEN_581;
  assign T_2723 = T_796 | T_1106;
  assign T_2724 = pageReplEn & T_2723;
  assign T_2726 = T_2724 != GEN_581;
  assign T_2727 = T_801 | T_1111;
  assign T_2728 = pageReplEn & T_2727;
  assign T_2730 = T_2728 != GEN_581;
  assign T_2731 = T_806 | T_1116;
  assign T_2732 = pageReplEn & T_2731;
  assign T_2734 = T_2732 != GEN_581;
  assign T_2735 = T_811 | T_1121;
  assign T_2736 = pageReplEn & T_2735;
  assign T_2738 = T_2736 != GEN_581;
  assign T_2739 = T_816 | T_1126;
  assign T_2740 = pageReplEn & T_2739;
  assign T_2742 = T_2740 != GEN_581;
  assign T_2743 = T_821 | T_1131;
  assign T_2744 = pageReplEn & T_2743;
  assign T_2746 = T_2744 != GEN_581;
  assign T_2747 = T_826 | T_1136;
  assign T_2748 = pageReplEn & T_2747;
  assign T_2750 = T_2748 != GEN_581;
  assign T_2751 = T_831 | T_1141;
  assign T_2752 = pageReplEn & T_2751;
  assign T_2754 = T_2752 != GEN_581;
  assign T_2755 = T_836 | T_1146;
  assign T_2756 = pageReplEn & T_2755;
  assign T_2758 = T_2756 != GEN_581;
  assign T_2759 = T_841 | T_1151;
  assign T_2760 = pageReplEn & T_2759;
  assign T_2762 = T_2760 != GEN_581;
  assign T_2763 = T_846 | T_1156;
  assign T_2764 = pageReplEn & T_2763;
  assign T_2766 = T_2764 != GEN_581;
  assign T_2767 = T_851 | T_1161;
  assign T_2768 = pageReplEn & T_2767;
  assign T_2770 = T_2768 != GEN_581;
  assign T_2771 = T_856 | T_1166;
  assign T_2772 = pageReplEn & T_2771;
  assign T_2774 = T_2772 != GEN_581;
  assign T_2775 = T_861 | T_1171;
  assign T_2776 = pageReplEn & T_2775;
  assign T_2778 = T_2776 != GEN_581;
  assign T_2779 = T_866 | T_1176;
  assign T_2780 = pageReplEn & T_2779;
  assign T_2782 = T_2780 != GEN_581;
  assign T_2783 = T_871 | T_1181;
  assign T_2784 = pageReplEn & T_2783;
  assign T_2786 = T_2784 != GEN_581;
  assign T_2787 = T_876 | T_1186;
  assign T_2788 = pageReplEn & T_2787;
  assign T_2790 = T_2788 != GEN_581;
  assign T_2791 = T_881 | T_1191;
  assign T_2792 = pageReplEn & T_2791;
  assign T_2794 = T_2792 != GEN_581;
  assign T_2795 = T_886 | T_1196;
  assign T_2796 = pageReplEn & T_2795;
  assign T_2798 = T_2796 != GEN_581;
  assign T_2804_0 = T_2554;
  assign T_2804_1 = T_2558;
  assign T_2804_2 = T_2562;
  assign T_2804_3 = T_2566;
  assign T_2804_4 = T_2570;
  assign T_2804_5 = T_2574;
  assign T_2804_6 = T_2578;
  assign T_2804_7 = T_2582;
  assign T_2804_8 = T_2586;
  assign T_2804_9 = T_2590;
  assign T_2804_10 = T_2594;
  assign T_2804_11 = T_2598;
  assign T_2804_12 = T_2602;
  assign T_2804_13 = T_2606;
  assign T_2804_14 = T_2610;
  assign T_2804_15 = T_2614;
  assign T_2804_16 = T_2618;
  assign T_2804_17 = T_2622;
  assign T_2804_18 = T_2626;
  assign T_2804_19 = T_2630;
  assign T_2804_20 = T_2634;
  assign T_2804_21 = T_2638;
  assign T_2804_22 = T_2642;
  assign T_2804_23 = T_2646;
  assign T_2804_24 = T_2650;
  assign T_2804_25 = T_2654;
  assign T_2804_26 = T_2658;
  assign T_2804_27 = T_2662;
  assign T_2804_28 = T_2666;
  assign T_2804_29 = T_2670;
  assign T_2804_30 = T_2674;
  assign T_2804_31 = T_2678;
  assign T_2804_32 = T_2682;
  assign T_2804_33 = T_2686;
  assign T_2804_34 = T_2690;
  assign T_2804_35 = T_2694;
  assign T_2804_36 = T_2698;
  assign T_2804_37 = T_2702;
  assign T_2804_38 = T_2706;
  assign T_2804_39 = T_2710;
  assign T_2804_40 = T_2714;
  assign T_2804_41 = T_2718;
  assign T_2804_42 = T_2722;
  assign T_2804_43 = T_2726;
  assign T_2804_44 = T_2730;
  assign T_2804_45 = T_2734;
  assign T_2804_46 = T_2738;
  assign T_2804_47 = T_2742;
  assign T_2804_48 = T_2746;
  assign T_2804_49 = T_2750;
  assign T_2804_50 = T_2754;
  assign T_2804_51 = T_2758;
  assign T_2804_52 = T_2762;
  assign T_2804_53 = T_2766;
  assign T_2804_54 = T_2770;
  assign T_2804_55 = T_2774;
  assign T_2804_56 = T_2778;
  assign T_2804_57 = T_2782;
  assign T_2804_58 = T_2786;
  assign T_2804_59 = T_2790;
  assign T_2804_60 = T_2794;
  assign T_2804_61 = T_2798;
  assign T_2806 = {T_2804_2,T_2804_1};
  assign T_2807 = {T_2806,T_2804_0};
  assign T_2808 = {T_2804_4,T_2804_3};
  assign T_2809 = {T_2804_6,T_2804_5};
  assign T_2810 = {T_2809,T_2808};
  assign T_2811 = {T_2810,T_2807};
  assign T_2812 = {T_2804_8,T_2804_7};
  assign T_2813 = {T_2804_10,T_2804_9};
  assign T_2814 = {T_2813,T_2812};
  assign T_2815 = {T_2804_12,T_2804_11};
  assign T_2816 = {T_2804_14,T_2804_13};
  assign T_2817 = {T_2816,T_2815};
  assign T_2818 = {T_2817,T_2814};
  assign T_2819 = {T_2818,T_2811};
  assign T_2820 = {T_2804_16,T_2804_15};
  assign T_2821 = {T_2804_18,T_2804_17};
  assign T_2822 = {T_2821,T_2820};
  assign T_2823 = {T_2804_20,T_2804_19};
  assign T_2824 = {T_2804_22,T_2804_21};
  assign T_2825 = {T_2824,T_2823};
  assign T_2826 = {T_2825,T_2822};
  assign T_2827 = {T_2804_24,T_2804_23};
  assign T_2828 = {T_2804_26,T_2804_25};
  assign T_2829 = {T_2828,T_2827};
  assign T_2830 = {T_2804_28,T_2804_27};
  assign T_2831 = {T_2804_30,T_2804_29};
  assign T_2832 = {T_2831,T_2830};
  assign T_2833 = {T_2832,T_2829};
  assign T_2834 = {T_2833,T_2826};
  assign T_2835 = {T_2834,T_2819};
  assign T_2836 = {T_2804_33,T_2804_32};
  assign T_2837 = {T_2836,T_2804_31};
  assign T_2838 = {T_2804_35,T_2804_34};
  assign T_2839 = {T_2804_37,T_2804_36};
  assign T_2840 = {T_2839,T_2838};
  assign T_2841 = {T_2840,T_2837};
  assign T_2842 = {T_2804_39,T_2804_38};
  assign T_2843 = {T_2804_41,T_2804_40};
  assign T_2844 = {T_2843,T_2842};
  assign T_2845 = {T_2804_43,T_2804_42};
  assign T_2846 = {T_2804_45,T_2804_44};
  assign T_2847 = {T_2846,T_2845};
  assign T_2848 = {T_2847,T_2844};
  assign T_2849 = {T_2848,T_2841};
  assign T_2850 = {T_2804_47,T_2804_46};
  assign T_2851 = {T_2804_49,T_2804_48};
  assign T_2852 = {T_2851,T_2850};
  assign T_2853 = {T_2804_51,T_2804_50};
  assign T_2854 = {T_2804_53,T_2804_52};
  assign T_2855 = {T_2854,T_2853};
  assign T_2856 = {T_2855,T_2852};
  assign T_2857 = {T_2804_55,T_2804_54};
  assign T_2858 = {T_2804_57,T_2804_56};
  assign T_2859 = {T_2858,T_2857};
  assign T_2860 = {T_2804_59,T_2804_58};
  assign T_2861 = {T_2804_61,T_2804_60};
  assign T_2862 = {T_2861,T_2860};
  assign T_2863 = {T_2862,T_2859};
  assign T_2864 = {T_2863,T_2856};
  assign T_2865 = {T_2864,T_2849};
  assign T_2866 = {T_2865,T_2835};
  assign GEN_780 = {{63'd0}, 1'h1};
  assign T_2868 = GEN_780 << T_2550;
  assign T_2869 = ~ T_2866;
  assign T_2870 = idxValid & T_2869;
  assign GEN_781 = {{2'd0}, T_2870};
  assign T_2871 = GEN_781 | T_2868;
  assign GEN_0 = r_btb_update_bits_isReturn;
  assign GEN_22 = GEN_581 == T_2550 ? GEN_0 : useRAS_0;
  assign GEN_23 = GEN_705 == T_2550 ? GEN_0 : useRAS_1;
  assign GEN_784 = {{4'd0}, 2'h2};
  assign GEN_24 = GEN_784 == T_2550 ? GEN_0 : useRAS_2;
  assign GEN_785 = {{4'd0}, 2'h3};
  assign GEN_25 = GEN_785 == T_2550 ? GEN_0 : useRAS_3;
  assign GEN_786 = {{3'd0}, 3'h4};
  assign GEN_26 = GEN_786 == T_2550 ? GEN_0 : useRAS_4;
  assign GEN_787 = {{3'd0}, 3'h5};
  assign GEN_27 = GEN_787 == T_2550 ? GEN_0 : useRAS_5;
  assign GEN_788 = {{3'd0}, 3'h6};
  assign GEN_28 = GEN_788 == T_2550 ? GEN_0 : useRAS_6;
  assign GEN_789 = {{3'd0}, 3'h7};
  assign GEN_29 = GEN_789 == T_2550 ? GEN_0 : useRAS_7;
  assign GEN_790 = {{2'd0}, 4'h8};
  assign GEN_30 = GEN_790 == T_2550 ? GEN_0 : useRAS_8;
  assign GEN_791 = {{2'd0}, 4'h9};
  assign GEN_31 = GEN_791 == T_2550 ? GEN_0 : useRAS_9;
  assign GEN_792 = {{2'd0}, 4'ha};
  assign GEN_32 = GEN_792 == T_2550 ? GEN_0 : useRAS_10;
  assign GEN_793 = {{2'd0}, 4'hb};
  assign GEN_33 = GEN_793 == T_2550 ? GEN_0 : useRAS_11;
  assign GEN_794 = {{2'd0}, 4'hc};
  assign GEN_34 = GEN_794 == T_2550 ? GEN_0 : useRAS_12;
  assign GEN_795 = {{2'd0}, 4'hd};
  assign GEN_35 = GEN_795 == T_2550 ? GEN_0 : useRAS_13;
  assign GEN_796 = {{2'd0}, 4'he};
  assign GEN_36 = GEN_796 == T_2550 ? GEN_0 : useRAS_14;
  assign GEN_797 = {{2'd0}, 4'hf};
  assign GEN_37 = GEN_797 == T_2550 ? GEN_0 : useRAS_15;
  assign GEN_798 = {{1'd0}, 5'h10};
  assign GEN_38 = GEN_798 == T_2550 ? GEN_0 : useRAS_16;
  assign GEN_799 = {{1'd0}, 5'h11};
  assign GEN_39 = GEN_799 == T_2550 ? GEN_0 : useRAS_17;
  assign GEN_800 = {{1'd0}, 5'h12};
  assign GEN_40 = GEN_800 == T_2550 ? GEN_0 : useRAS_18;
  assign GEN_801 = {{1'd0}, 5'h13};
  assign GEN_41 = GEN_801 == T_2550 ? GEN_0 : useRAS_19;
  assign GEN_802 = {{1'd0}, 5'h14};
  assign GEN_42 = GEN_802 == T_2550 ? GEN_0 : useRAS_20;
  assign GEN_803 = {{1'd0}, 5'h15};
  assign GEN_43 = GEN_803 == T_2550 ? GEN_0 : useRAS_21;
  assign GEN_804 = {{1'd0}, 5'h16};
  assign GEN_44 = GEN_804 == T_2550 ? GEN_0 : useRAS_22;
  assign GEN_805 = {{1'd0}, 5'h17};
  assign GEN_45 = GEN_805 == T_2550 ? GEN_0 : useRAS_23;
  assign GEN_806 = {{1'd0}, 5'h18};
  assign GEN_46 = GEN_806 == T_2550 ? GEN_0 : useRAS_24;
  assign GEN_807 = {{1'd0}, 5'h19};
  assign GEN_47 = GEN_807 == T_2550 ? GEN_0 : useRAS_25;
  assign GEN_808 = {{1'd0}, 5'h1a};
  assign GEN_48 = GEN_808 == T_2550 ? GEN_0 : useRAS_26;
  assign GEN_809 = {{1'd0}, 5'h1b};
  assign GEN_49 = GEN_809 == T_2550 ? GEN_0 : useRAS_27;
  assign GEN_810 = {{1'd0}, 5'h1c};
  assign GEN_50 = GEN_810 == T_2550 ? GEN_0 : useRAS_28;
  assign GEN_811 = {{1'd0}, 5'h1d};
  assign GEN_51 = GEN_811 == T_2550 ? GEN_0 : useRAS_29;
  assign GEN_812 = {{1'd0}, 5'h1e};
  assign GEN_52 = GEN_812 == T_2550 ? GEN_0 : useRAS_30;
  assign GEN_813 = {{1'd0}, 5'h1f};
  assign GEN_53 = GEN_813 == T_2550 ? GEN_0 : useRAS_31;
  assign GEN_54 = 6'h20 == T_2550 ? GEN_0 : useRAS_32;
  assign GEN_55 = 6'h21 == T_2550 ? GEN_0 : useRAS_33;
  assign GEN_56 = 6'h22 == T_2550 ? GEN_0 : useRAS_34;
  assign GEN_57 = 6'h23 == T_2550 ? GEN_0 : useRAS_35;
  assign GEN_58 = 6'h24 == T_2550 ? GEN_0 : useRAS_36;
  assign GEN_59 = 6'h25 == T_2550 ? GEN_0 : useRAS_37;
  assign GEN_60 = 6'h26 == T_2550 ? GEN_0 : useRAS_38;
  assign GEN_61 = 6'h27 == T_2550 ? GEN_0 : useRAS_39;
  assign GEN_62 = 6'h28 == T_2550 ? GEN_0 : useRAS_40;
  assign GEN_63 = 6'h29 == T_2550 ? GEN_0 : useRAS_41;
  assign GEN_64 = 6'h2a == T_2550 ? GEN_0 : useRAS_42;
  assign GEN_65 = 6'h2b == T_2550 ? GEN_0 : useRAS_43;
  assign GEN_66 = 6'h2c == T_2550 ? GEN_0 : useRAS_44;
  assign GEN_67 = 6'h2d == T_2550 ? GEN_0 : useRAS_45;
  assign GEN_68 = 6'h2e == T_2550 ? GEN_0 : useRAS_46;
  assign GEN_69 = 6'h2f == T_2550 ? GEN_0 : useRAS_47;
  assign GEN_70 = 6'h30 == T_2550 ? GEN_0 : useRAS_48;
  assign GEN_71 = 6'h31 == T_2550 ? GEN_0 : useRAS_49;
  assign GEN_72 = 6'h32 == T_2550 ? GEN_0 : useRAS_50;
  assign GEN_73 = 6'h33 == T_2550 ? GEN_0 : useRAS_51;
  assign GEN_74 = 6'h34 == T_2550 ? GEN_0 : useRAS_52;
  assign GEN_75 = 6'h35 == T_2550 ? GEN_0 : useRAS_53;
  assign GEN_76 = 6'h36 == T_2550 ? GEN_0 : useRAS_54;
  assign GEN_77 = 6'h37 == T_2550 ? GEN_0 : useRAS_55;
  assign GEN_78 = 6'h38 == T_2550 ? GEN_0 : useRAS_56;
  assign GEN_79 = 6'h39 == T_2550 ? GEN_0 : useRAS_57;
  assign GEN_80 = 6'h3a == T_2550 ? GEN_0 : useRAS_58;
  assign GEN_81 = 6'h3b == T_2550 ? GEN_0 : useRAS_59;
  assign GEN_82 = 6'h3c == T_2550 ? GEN_0 : useRAS_60;
  assign GEN_83 = 6'h3d == T_2550 ? GEN_0 : useRAS_61;
  assign GEN_1 = r_btb_update_bits_isJump;
  assign GEN_84 = GEN_581 == T_2550 ? GEN_1 : isJump_0;
  assign GEN_85 = GEN_705 == T_2550 ? GEN_1 : isJump_1;
  assign GEN_86 = GEN_784 == T_2550 ? GEN_1 : isJump_2;
  assign GEN_87 = GEN_785 == T_2550 ? GEN_1 : isJump_3;
  assign GEN_88 = GEN_786 == T_2550 ? GEN_1 : isJump_4;
  assign GEN_89 = GEN_787 == T_2550 ? GEN_1 : isJump_5;
  assign GEN_90 = GEN_788 == T_2550 ? GEN_1 : isJump_6;
  assign GEN_91 = GEN_789 == T_2550 ? GEN_1 : isJump_7;
  assign GEN_92 = GEN_790 == T_2550 ? GEN_1 : isJump_8;
  assign GEN_93 = GEN_791 == T_2550 ? GEN_1 : isJump_9;
  assign GEN_94 = GEN_792 == T_2550 ? GEN_1 : isJump_10;
  assign GEN_95 = GEN_793 == T_2550 ? GEN_1 : isJump_11;
  assign GEN_96 = GEN_794 == T_2550 ? GEN_1 : isJump_12;
  assign GEN_97 = GEN_795 == T_2550 ? GEN_1 : isJump_13;
  assign GEN_98 = GEN_796 == T_2550 ? GEN_1 : isJump_14;
  assign GEN_99 = GEN_797 == T_2550 ? GEN_1 : isJump_15;
  assign GEN_100 = GEN_798 == T_2550 ? GEN_1 : isJump_16;
  assign GEN_101 = GEN_799 == T_2550 ? GEN_1 : isJump_17;
  assign GEN_102 = GEN_800 == T_2550 ? GEN_1 : isJump_18;
  assign GEN_103 = GEN_801 == T_2550 ? GEN_1 : isJump_19;
  assign GEN_104 = GEN_802 == T_2550 ? GEN_1 : isJump_20;
  assign GEN_105 = GEN_803 == T_2550 ? GEN_1 : isJump_21;
  assign GEN_106 = GEN_804 == T_2550 ? GEN_1 : isJump_22;
  assign GEN_107 = GEN_805 == T_2550 ? GEN_1 : isJump_23;
  assign GEN_108 = GEN_806 == T_2550 ? GEN_1 : isJump_24;
  assign GEN_109 = GEN_807 == T_2550 ? GEN_1 : isJump_25;
  assign GEN_110 = GEN_808 == T_2550 ? GEN_1 : isJump_26;
  assign GEN_111 = GEN_809 == T_2550 ? GEN_1 : isJump_27;
  assign GEN_112 = GEN_810 == T_2550 ? GEN_1 : isJump_28;
  assign GEN_113 = GEN_811 == T_2550 ? GEN_1 : isJump_29;
  assign GEN_114 = GEN_812 == T_2550 ? GEN_1 : isJump_30;
  assign GEN_115 = GEN_813 == T_2550 ? GEN_1 : isJump_31;
  assign GEN_116 = 6'h20 == T_2550 ? GEN_1 : isJump_32;
  assign GEN_117 = 6'h21 == T_2550 ? GEN_1 : isJump_33;
  assign GEN_118 = 6'h22 == T_2550 ? GEN_1 : isJump_34;
  assign GEN_119 = 6'h23 == T_2550 ? GEN_1 : isJump_35;
  assign GEN_120 = 6'h24 == T_2550 ? GEN_1 : isJump_36;
  assign GEN_121 = 6'h25 == T_2550 ? GEN_1 : isJump_37;
  assign GEN_122 = 6'h26 == T_2550 ? GEN_1 : isJump_38;
  assign GEN_123 = 6'h27 == T_2550 ? GEN_1 : isJump_39;
  assign GEN_124 = 6'h28 == T_2550 ? GEN_1 : isJump_40;
  assign GEN_125 = 6'h29 == T_2550 ? GEN_1 : isJump_41;
  assign GEN_126 = 6'h2a == T_2550 ? GEN_1 : isJump_42;
  assign GEN_127 = 6'h2b == T_2550 ? GEN_1 : isJump_43;
  assign GEN_128 = 6'h2c == T_2550 ? GEN_1 : isJump_44;
  assign GEN_129 = 6'h2d == T_2550 ? GEN_1 : isJump_45;
  assign GEN_130 = 6'h2e == T_2550 ? GEN_1 : isJump_46;
  assign GEN_131 = 6'h2f == T_2550 ? GEN_1 : isJump_47;
  assign GEN_132 = 6'h30 == T_2550 ? GEN_1 : isJump_48;
  assign GEN_133 = 6'h31 == T_2550 ? GEN_1 : isJump_49;
  assign GEN_134 = 6'h32 == T_2550 ? GEN_1 : isJump_50;
  assign GEN_135 = 6'h33 == T_2550 ? GEN_1 : isJump_51;
  assign GEN_136 = 6'h34 == T_2550 ? GEN_1 : isJump_52;
  assign GEN_137 = 6'h35 == T_2550 ? GEN_1 : isJump_53;
  assign GEN_138 = 6'h36 == T_2550 ? GEN_1 : isJump_54;
  assign GEN_139 = 6'h37 == T_2550 ? GEN_1 : isJump_55;
  assign GEN_140 = 6'h38 == T_2550 ? GEN_1 : isJump_56;
  assign GEN_141 = 6'h39 == T_2550 ? GEN_1 : isJump_57;
  assign GEN_142 = 6'h3a == T_2550 ? GEN_1 : isJump_58;
  assign GEN_143 = 6'h3b == T_2550 ? GEN_1 : isJump_59;
  assign GEN_144 = 6'h3c == T_2550 ? GEN_1 : isJump_60;
  assign GEN_145 = 6'h3d == T_2550 ? GEN_1 : isJump_61;
  assign T_2881 = idxPageUpdateOH & 6'h15;
  assign T_2883 = T_2881 != GEN_581;
  assign T_2884 = T_2883 ? doIdxPageRepl : doTgtPageRepl;
  assign T_2887 = T_2883 ? T_1939 : T_1398;
  assign T_2888 = pageReplEn[0];
  assign T_2889 = T_2884 & T_2888;
  assign T_2892 = pageReplEn[2];
  assign T_2893 = T_2884 & T_2892;
  assign T_2896 = pageReplEn[4];
  assign T_2897 = T_2884 & T_2896;
  assign T_2900 = T_2883 ? doTgtPageRepl : doIdxPageRepl;
  assign T_2903 = T_2883 ? T_1398 : T_1939;
  assign T_2904 = pageReplEn[1];
  assign T_2905 = T_2900 & T_2904;
  assign T_2908 = pageReplEn[3];
  assign T_2909 = T_2900 & T_2908;
  assign T_2912 = pageReplEn[5];
  assign T_2913 = T_2900 & T_2912;
  assign T_2916 = pageValid | pageReplEn;
  assign GEN_176 = doPageRepl ? T_2916 : pageValid;
  assign GEN_239 = r_btb_update_valid ? T_2871 : {{2'd0}, idxValid};
  assign GEN_261 = r_btb_update_valid ? GEN_22 : useRAS_0;
  assign GEN_262 = r_btb_update_valid ? GEN_23 : useRAS_1;
  assign GEN_263 = r_btb_update_valid ? GEN_24 : useRAS_2;
  assign GEN_264 = r_btb_update_valid ? GEN_25 : useRAS_3;
  assign GEN_265 = r_btb_update_valid ? GEN_26 : useRAS_4;
  assign GEN_266 = r_btb_update_valid ? GEN_27 : useRAS_5;
  assign GEN_267 = r_btb_update_valid ? GEN_28 : useRAS_6;
  assign GEN_268 = r_btb_update_valid ? GEN_29 : useRAS_7;
  assign GEN_269 = r_btb_update_valid ? GEN_30 : useRAS_8;
  assign GEN_270 = r_btb_update_valid ? GEN_31 : useRAS_9;
  assign GEN_271 = r_btb_update_valid ? GEN_32 : useRAS_10;
  assign GEN_272 = r_btb_update_valid ? GEN_33 : useRAS_11;
  assign GEN_273 = r_btb_update_valid ? GEN_34 : useRAS_12;
  assign GEN_274 = r_btb_update_valid ? GEN_35 : useRAS_13;
  assign GEN_275 = r_btb_update_valid ? GEN_36 : useRAS_14;
  assign GEN_276 = r_btb_update_valid ? GEN_37 : useRAS_15;
  assign GEN_277 = r_btb_update_valid ? GEN_38 : useRAS_16;
  assign GEN_278 = r_btb_update_valid ? GEN_39 : useRAS_17;
  assign GEN_279 = r_btb_update_valid ? GEN_40 : useRAS_18;
  assign GEN_280 = r_btb_update_valid ? GEN_41 : useRAS_19;
  assign GEN_281 = r_btb_update_valid ? GEN_42 : useRAS_20;
  assign GEN_282 = r_btb_update_valid ? GEN_43 : useRAS_21;
  assign GEN_283 = r_btb_update_valid ? GEN_44 : useRAS_22;
  assign GEN_284 = r_btb_update_valid ? GEN_45 : useRAS_23;
  assign GEN_285 = r_btb_update_valid ? GEN_46 : useRAS_24;
  assign GEN_286 = r_btb_update_valid ? GEN_47 : useRAS_25;
  assign GEN_287 = r_btb_update_valid ? GEN_48 : useRAS_26;
  assign GEN_288 = r_btb_update_valid ? GEN_49 : useRAS_27;
  assign GEN_289 = r_btb_update_valid ? GEN_50 : useRAS_28;
  assign GEN_290 = r_btb_update_valid ? GEN_51 : useRAS_29;
  assign GEN_291 = r_btb_update_valid ? GEN_52 : useRAS_30;
  assign GEN_292 = r_btb_update_valid ? GEN_53 : useRAS_31;
  assign GEN_293 = r_btb_update_valid ? GEN_54 : useRAS_32;
  assign GEN_294 = r_btb_update_valid ? GEN_55 : useRAS_33;
  assign GEN_295 = r_btb_update_valid ? GEN_56 : useRAS_34;
  assign GEN_296 = r_btb_update_valid ? GEN_57 : useRAS_35;
  assign GEN_297 = r_btb_update_valid ? GEN_58 : useRAS_36;
  assign GEN_298 = r_btb_update_valid ? GEN_59 : useRAS_37;
  assign GEN_299 = r_btb_update_valid ? GEN_60 : useRAS_38;
  assign GEN_300 = r_btb_update_valid ? GEN_61 : useRAS_39;
  assign GEN_301 = r_btb_update_valid ? GEN_62 : useRAS_40;
  assign GEN_302 = r_btb_update_valid ? GEN_63 : useRAS_41;
  assign GEN_303 = r_btb_update_valid ? GEN_64 : useRAS_42;
  assign GEN_304 = r_btb_update_valid ? GEN_65 : useRAS_43;
  assign GEN_305 = r_btb_update_valid ? GEN_66 : useRAS_44;
  assign GEN_306 = r_btb_update_valid ? GEN_67 : useRAS_45;
  assign GEN_307 = r_btb_update_valid ? GEN_68 : useRAS_46;
  assign GEN_308 = r_btb_update_valid ? GEN_69 : useRAS_47;
  assign GEN_309 = r_btb_update_valid ? GEN_70 : useRAS_48;
  assign GEN_310 = r_btb_update_valid ? GEN_71 : useRAS_49;
  assign GEN_311 = r_btb_update_valid ? GEN_72 : useRAS_50;
  assign GEN_312 = r_btb_update_valid ? GEN_73 : useRAS_51;
  assign GEN_313 = r_btb_update_valid ? GEN_74 : useRAS_52;
  assign GEN_314 = r_btb_update_valid ? GEN_75 : useRAS_53;
  assign GEN_315 = r_btb_update_valid ? GEN_76 : useRAS_54;
  assign GEN_316 = r_btb_update_valid ? GEN_77 : useRAS_55;
  assign GEN_317 = r_btb_update_valid ? GEN_78 : useRAS_56;
  assign GEN_318 = r_btb_update_valid ? GEN_79 : useRAS_57;
  assign GEN_319 = r_btb_update_valid ? GEN_80 : useRAS_58;
  assign GEN_320 = r_btb_update_valid ? GEN_81 : useRAS_59;
  assign GEN_321 = r_btb_update_valid ? GEN_82 : useRAS_60;
  assign GEN_322 = r_btb_update_valid ? GEN_83 : useRAS_61;
  assign GEN_324 = r_btb_update_valid ? GEN_84 : isJump_0;
  assign GEN_325 = r_btb_update_valid ? GEN_85 : isJump_1;
  assign GEN_326 = r_btb_update_valid ? GEN_86 : isJump_2;
  assign GEN_327 = r_btb_update_valid ? GEN_87 : isJump_3;
  assign GEN_328 = r_btb_update_valid ? GEN_88 : isJump_4;
  assign GEN_329 = r_btb_update_valid ? GEN_89 : isJump_5;
  assign GEN_330 = r_btb_update_valid ? GEN_90 : isJump_6;
  assign GEN_331 = r_btb_update_valid ? GEN_91 : isJump_7;
  assign GEN_332 = r_btb_update_valid ? GEN_92 : isJump_8;
  assign GEN_333 = r_btb_update_valid ? GEN_93 : isJump_9;
  assign GEN_334 = r_btb_update_valid ? GEN_94 : isJump_10;
  assign GEN_335 = r_btb_update_valid ? GEN_95 : isJump_11;
  assign GEN_336 = r_btb_update_valid ? GEN_96 : isJump_12;
  assign GEN_337 = r_btb_update_valid ? GEN_97 : isJump_13;
  assign GEN_338 = r_btb_update_valid ? GEN_98 : isJump_14;
  assign GEN_339 = r_btb_update_valid ? GEN_99 : isJump_15;
  assign GEN_340 = r_btb_update_valid ? GEN_100 : isJump_16;
  assign GEN_341 = r_btb_update_valid ? GEN_101 : isJump_17;
  assign GEN_342 = r_btb_update_valid ? GEN_102 : isJump_18;
  assign GEN_343 = r_btb_update_valid ? GEN_103 : isJump_19;
  assign GEN_344 = r_btb_update_valid ? GEN_104 : isJump_20;
  assign GEN_345 = r_btb_update_valid ? GEN_105 : isJump_21;
  assign GEN_346 = r_btb_update_valid ? GEN_106 : isJump_22;
  assign GEN_347 = r_btb_update_valid ? GEN_107 : isJump_23;
  assign GEN_348 = r_btb_update_valid ? GEN_108 : isJump_24;
  assign GEN_349 = r_btb_update_valid ? GEN_109 : isJump_25;
  assign GEN_350 = r_btb_update_valid ? GEN_110 : isJump_26;
  assign GEN_351 = r_btb_update_valid ? GEN_111 : isJump_27;
  assign GEN_352 = r_btb_update_valid ? GEN_112 : isJump_28;
  assign GEN_353 = r_btb_update_valid ? GEN_113 : isJump_29;
  assign GEN_354 = r_btb_update_valid ? GEN_114 : isJump_30;
  assign GEN_355 = r_btb_update_valid ? GEN_115 : isJump_31;
  assign GEN_356 = r_btb_update_valid ? GEN_116 : isJump_32;
  assign GEN_357 = r_btb_update_valid ? GEN_117 : isJump_33;
  assign GEN_358 = r_btb_update_valid ? GEN_118 : isJump_34;
  assign GEN_359 = r_btb_update_valid ? GEN_119 : isJump_35;
  assign GEN_360 = r_btb_update_valid ? GEN_120 : isJump_36;
  assign GEN_361 = r_btb_update_valid ? GEN_121 : isJump_37;
  assign GEN_362 = r_btb_update_valid ? GEN_122 : isJump_38;
  assign GEN_363 = r_btb_update_valid ? GEN_123 : isJump_39;
  assign GEN_364 = r_btb_update_valid ? GEN_124 : isJump_40;
  assign GEN_365 = r_btb_update_valid ? GEN_125 : isJump_41;
  assign GEN_366 = r_btb_update_valid ? GEN_126 : isJump_42;
  assign GEN_367 = r_btb_update_valid ? GEN_127 : isJump_43;
  assign GEN_368 = r_btb_update_valid ? GEN_128 : isJump_44;
  assign GEN_369 = r_btb_update_valid ? GEN_129 : isJump_45;
  assign GEN_370 = r_btb_update_valid ? GEN_130 : isJump_46;
  assign GEN_371 = r_btb_update_valid ? GEN_131 : isJump_47;
  assign GEN_372 = r_btb_update_valid ? GEN_132 : isJump_48;
  assign GEN_373 = r_btb_update_valid ? GEN_133 : isJump_49;
  assign GEN_374 = r_btb_update_valid ? GEN_134 : isJump_50;
  assign GEN_375 = r_btb_update_valid ? GEN_135 : isJump_51;
  assign GEN_376 = r_btb_update_valid ? GEN_136 : isJump_52;
  assign GEN_377 = r_btb_update_valid ? GEN_137 : isJump_53;
  assign GEN_378 = r_btb_update_valid ? GEN_138 : isJump_54;
  assign GEN_379 = r_btb_update_valid ? GEN_139 : isJump_55;
  assign GEN_380 = r_btb_update_valid ? GEN_140 : isJump_56;
  assign GEN_381 = r_btb_update_valid ? GEN_141 : isJump_57;
  assign GEN_382 = r_btb_update_valid ? GEN_142 : isJump_58;
  assign GEN_383 = r_btb_update_valid ? GEN_143 : isJump_59;
  assign GEN_384 = r_btb_update_valid ? GEN_144 : isJump_60;
  assign GEN_385 = r_btb_update_valid ? GEN_145 : isJump_61;
  assign GEN_393 = r_btb_update_valid ? T_2889 : 1'h0;
  assign GEN_398 = r_btb_update_valid ? T_2893 : 1'h0;
  assign GEN_403 = r_btb_update_valid ? T_2897 : 1'h0;
  assign GEN_408 = r_btb_update_valid ? T_2905 : 1'h0;
  assign GEN_413 = r_btb_update_valid ? T_2909 : 1'h0;
  assign GEN_418 = r_btb_update_valid ? T_2913 : 1'h0;
  assign GEN_421 = r_btb_update_valid ? GEN_176 : pageValid;
  assign GEN_422 = io_invalidate ? {{63'd0}, 1'h0} : GEN_239;
  assign GEN_423 = io_invalidate ? {{5'd0}, 1'h0} : GEN_421;
  assign GEN_847 = {{61'd0}, 1'h0};
  assign T_2920 = hits != GEN_847;
  assign T_2921 = hits[0];
  assign T_2922 = hits[1];
  assign T_2923 = hits[2];
  assign T_2924 = hits[3];
  assign T_2925 = hits[4];
  assign T_2926 = hits[5];
  assign T_2927 = hits[6];
  assign T_2928 = hits[7];
  assign T_2929 = hits[8];
  assign T_2930 = hits[9];
  assign T_2931 = hits[10];
  assign T_2932 = hits[11];
  assign T_2933 = hits[12];
  assign T_2934 = hits[13];
  assign T_2935 = hits[14];
  assign T_2936 = hits[15];
  assign T_2937 = hits[16];
  assign T_2938 = hits[17];
  assign T_2939 = hits[18];
  assign T_2940 = hits[19];
  assign T_2941 = hits[20];
  assign T_2942 = hits[21];
  assign T_2943 = hits[22];
  assign T_2944 = hits[23];
  assign T_2945 = hits[24];
  assign T_2946 = hits[25];
  assign T_2947 = hits[26];
  assign T_2948 = hits[27];
  assign T_2949 = hits[28];
  assign T_2950 = hits[29];
  assign T_2951 = hits[30];
  assign T_2952 = hits[31];
  assign T_2953 = hits[32];
  assign T_2954 = hits[33];
  assign T_2955 = hits[34];
  assign T_2956 = hits[35];
  assign T_2957 = hits[36];
  assign T_2958 = hits[37];
  assign T_2959 = hits[38];
  assign T_2960 = hits[39];
  assign T_2961 = hits[40];
  assign T_2962 = hits[41];
  assign T_2963 = hits[42];
  assign T_2964 = hits[43];
  assign T_2965 = hits[44];
  assign T_2966 = hits[45];
  assign T_2967 = hits[46];
  assign T_2968 = hits[47];
  assign T_2969 = hits[48];
  assign T_2970 = hits[49];
  assign T_2971 = hits[50];
  assign T_2972 = hits[51];
  assign T_2973 = hits[52];
  assign T_2974 = hits[53];
  assign T_2975 = hits[54];
  assign T_2976 = hits[55];
  assign T_2977 = hits[56];
  assign T_2978 = hits[57];
  assign T_2979 = hits[58];
  assign T_2980 = hits[59];
  assign T_2981 = hits[60];
  assign T_2982 = hits[61];
  assign T_2984 = T_2921 ? T_891 : {{5'd0}, 1'h0};
  assign T_2986 = T_2922 ? T_896 : {{5'd0}, 1'h0};
  assign T_2988 = T_2923 ? T_901 : {{5'd0}, 1'h0};
  assign T_2990 = T_2924 ? T_906 : {{5'd0}, 1'h0};
  assign T_2992 = T_2925 ? T_911 : {{5'd0}, 1'h0};
  assign T_2994 = T_2926 ? T_916 : {{5'd0}, 1'h0};
  assign T_2996 = T_2927 ? T_921 : {{5'd0}, 1'h0};
  assign T_2998 = T_2928 ? T_926 : {{5'd0}, 1'h0};
  assign T_3000 = T_2929 ? T_931 : {{5'd0}, 1'h0};
  assign T_3002 = T_2930 ? T_936 : {{5'd0}, 1'h0};
  assign T_3004 = T_2931 ? T_941 : {{5'd0}, 1'h0};
  assign T_3006 = T_2932 ? T_946 : {{5'd0}, 1'h0};
  assign T_3008 = T_2933 ? T_951 : {{5'd0}, 1'h0};
  assign T_3010 = T_2934 ? T_956 : {{5'd0}, 1'h0};
  assign T_3012 = T_2935 ? T_961 : {{5'd0}, 1'h0};
  assign T_3014 = T_2936 ? T_966 : {{5'd0}, 1'h0};
  assign T_3016 = T_2937 ? T_971 : {{5'd0}, 1'h0};
  assign T_3018 = T_2938 ? T_976 : {{5'd0}, 1'h0};
  assign T_3020 = T_2939 ? T_981 : {{5'd0}, 1'h0};
  assign T_3022 = T_2940 ? T_986 : {{5'd0}, 1'h0};
  assign T_3024 = T_2941 ? T_991 : {{5'd0}, 1'h0};
  assign T_3026 = T_2942 ? T_996 : {{5'd0}, 1'h0};
  assign T_3028 = T_2943 ? T_1001 : {{5'd0}, 1'h0};
  assign T_3030 = T_2944 ? T_1006 : {{5'd0}, 1'h0};
  assign T_3032 = T_2945 ? T_1011 : {{5'd0}, 1'h0};
  assign T_3034 = T_2946 ? T_1016 : {{5'd0}, 1'h0};
  assign T_3036 = T_2947 ? T_1021 : {{5'd0}, 1'h0};
  assign T_3038 = T_2948 ? T_1026 : {{5'd0}, 1'h0};
  assign T_3040 = T_2949 ? T_1031 : {{5'd0}, 1'h0};
  assign T_3042 = T_2950 ? T_1036 : {{5'd0}, 1'h0};
  assign T_3044 = T_2951 ? T_1041 : {{5'd0}, 1'h0};
  assign T_3046 = T_2952 ? T_1046 : {{5'd0}, 1'h0};
  assign T_3048 = T_2953 ? T_1051 : {{5'd0}, 1'h0};
  assign T_3050 = T_2954 ? T_1056 : {{5'd0}, 1'h0};
  assign T_3052 = T_2955 ? T_1061 : {{5'd0}, 1'h0};
  assign T_3054 = T_2956 ? T_1066 : {{5'd0}, 1'h0};
  assign T_3056 = T_2957 ? T_1071 : {{5'd0}, 1'h0};
  assign T_3058 = T_2958 ? T_1076 : {{5'd0}, 1'h0};
  assign T_3060 = T_2959 ? T_1081 : {{5'd0}, 1'h0};
  assign T_3062 = T_2960 ? T_1086 : {{5'd0}, 1'h0};
  assign T_3064 = T_2961 ? T_1091 : {{5'd0}, 1'h0};
  assign T_3066 = T_2962 ? T_1096 : {{5'd0}, 1'h0};
  assign T_3068 = T_2963 ? T_1101 : {{5'd0}, 1'h0};
  assign T_3070 = T_2964 ? T_1106 : {{5'd0}, 1'h0};
  assign T_3072 = T_2965 ? T_1111 : {{5'd0}, 1'h0};
  assign T_3074 = T_2966 ? T_1116 : {{5'd0}, 1'h0};
  assign T_3076 = T_2967 ? T_1121 : {{5'd0}, 1'h0};
  assign T_3078 = T_2968 ? T_1126 : {{5'd0}, 1'h0};
  assign T_3080 = T_2969 ? T_1131 : {{5'd0}, 1'h0};
  assign T_3082 = T_2970 ? T_1136 : {{5'd0}, 1'h0};
  assign T_3084 = T_2971 ? T_1141 : {{5'd0}, 1'h0};
  assign T_3086 = T_2972 ? T_1146 : {{5'd0}, 1'h0};
  assign T_3088 = T_2973 ? T_1151 : {{5'd0}, 1'h0};
  assign T_3090 = T_2974 ? T_1156 : {{5'd0}, 1'h0};
  assign T_3092 = T_2975 ? T_1161 : {{5'd0}, 1'h0};
  assign T_3094 = T_2976 ? T_1166 : {{5'd0}, 1'h0};
  assign T_3096 = T_2977 ? T_1171 : {{5'd0}, 1'h0};
  assign T_3098 = T_2978 ? T_1176 : {{5'd0}, 1'h0};
  assign T_3100 = T_2979 ? T_1181 : {{5'd0}, 1'h0};
  assign T_3102 = T_2980 ? T_1186 : {{5'd0}, 1'h0};
  assign T_3104 = T_2981 ? T_1191 : {{5'd0}, 1'h0};
  assign T_3106 = T_2982 ? T_1196 : {{5'd0}, 1'h0};
  assign T_3108 = T_2984 | T_2986;
  assign T_3109 = T_3108 | T_2988;
  assign T_3110 = T_3109 | T_2990;
  assign T_3111 = T_3110 | T_2992;
  assign T_3112 = T_3111 | T_2994;
  assign T_3113 = T_3112 | T_2996;
  assign T_3114 = T_3113 | T_2998;
  assign T_3115 = T_3114 | T_3000;
  assign T_3116 = T_3115 | T_3002;
  assign T_3117 = T_3116 | T_3004;
  assign T_3118 = T_3117 | T_3006;
  assign T_3119 = T_3118 | T_3008;
  assign T_3120 = T_3119 | T_3010;
  assign T_3121 = T_3120 | T_3012;
  assign T_3122 = T_3121 | T_3014;
  assign T_3123 = T_3122 | T_3016;
  assign T_3124 = T_3123 | T_3018;
  assign T_3125 = T_3124 | T_3020;
  assign T_3126 = T_3125 | T_3022;
  assign T_3127 = T_3126 | T_3024;
  assign T_3128 = T_3127 | T_3026;
  assign T_3129 = T_3128 | T_3028;
  assign T_3130 = T_3129 | T_3030;
  assign T_3131 = T_3130 | T_3032;
  assign T_3132 = T_3131 | T_3034;
  assign T_3133 = T_3132 | T_3036;
  assign T_3134 = T_3133 | T_3038;
  assign T_3135 = T_3134 | T_3040;
  assign T_3136 = T_3135 | T_3042;
  assign T_3137 = T_3136 | T_3044;
  assign T_3138 = T_3137 | T_3046;
  assign T_3139 = T_3138 | T_3048;
  assign T_3140 = T_3139 | T_3050;
  assign T_3141 = T_3140 | T_3052;
  assign T_3142 = T_3141 | T_3054;
  assign T_3143 = T_3142 | T_3056;
  assign T_3144 = T_3143 | T_3058;
  assign T_3145 = T_3144 | T_3060;
  assign T_3146 = T_3145 | T_3062;
  assign T_3147 = T_3146 | T_3064;
  assign T_3148 = T_3147 | T_3066;
  assign T_3149 = T_3148 | T_3068;
  assign T_3150 = T_3149 | T_3070;
  assign T_3151 = T_3150 | T_3072;
  assign T_3152 = T_3151 | T_3074;
  assign T_3153 = T_3152 | T_3076;
  assign T_3154 = T_3153 | T_3078;
  assign T_3155 = T_3154 | T_3080;
  assign T_3156 = T_3155 | T_3082;
  assign T_3157 = T_3156 | T_3084;
  assign T_3158 = T_3157 | T_3086;
  assign T_3159 = T_3158 | T_3088;
  assign T_3160 = T_3159 | T_3090;
  assign T_3161 = T_3160 | T_3092;
  assign T_3162 = T_3161 | T_3094;
  assign T_3163 = T_3162 | T_3096;
  assign T_3164 = T_3163 | T_3098;
  assign T_3165 = T_3164 | T_3100;
  assign T_3166 = T_3165 | T_3102;
  assign T_3167 = T_3166 | T_3104;
  assign T_3168 = T_3167 | T_3106;
  assign T_3169 = T_3168;
  assign T_3170 = T_3169[0];
  assign T_3171 = T_3169[1];
  assign T_3172 = T_3169[2];
  assign T_3173 = T_3169[3];
  assign T_3174 = T_3169[4];
  assign T_3175 = T_3169[5];
  assign T_3189 = T_3170 ? pages_T_3177_data : {{26'd0}, 1'h0};
  assign T_3191 = T_3171 ? pages_T_3179_data : {{26'd0}, 1'h0};
  assign T_3193 = T_3172 ? pages_T_3181_data : {{26'd0}, 1'h0};
  assign T_3195 = T_3173 ? pages_T_3183_data : {{26'd0}, 1'h0};
  assign T_3197 = T_3174 ? pages_T_3185_data : {{26'd0}, 1'h0};
  assign T_3199 = T_3175 ? pages_T_3187_data : {{26'd0}, 1'h0};
  assign T_3201 = T_3189 | T_3191;
  assign T_3202 = T_3201 | T_3193;
  assign T_3203 = T_3202 | T_3195;
  assign T_3204 = T_3203 | T_3197;
  assign T_3205 = T_3204 | T_3199;
  assign T_3206 = T_3205;
  assign T_3394 = T_2921 ? tgts_T_3270_data : {{11'd0}, 1'h0};
  assign T_3396 = T_2922 ? tgts_T_3272_data : {{11'd0}, 1'h0};
  assign T_3398 = T_2923 ? tgts_T_3274_data : {{11'd0}, 1'h0};
  assign T_3400 = T_2924 ? tgts_T_3276_data : {{11'd0}, 1'h0};
  assign T_3402 = T_2925 ? tgts_T_3278_data : {{11'd0}, 1'h0};
  assign T_3404 = T_2926 ? tgts_T_3280_data : {{11'd0}, 1'h0};
  assign T_3406 = T_2927 ? tgts_T_3282_data : {{11'd0}, 1'h0};
  assign T_3408 = T_2928 ? tgts_T_3284_data : {{11'd0}, 1'h0};
  assign T_3410 = T_2929 ? tgts_T_3286_data : {{11'd0}, 1'h0};
  assign T_3412 = T_2930 ? tgts_T_3288_data : {{11'd0}, 1'h0};
  assign T_3414 = T_2931 ? tgts_T_3290_data : {{11'd0}, 1'h0};
  assign T_3416 = T_2932 ? tgts_T_3292_data : {{11'd0}, 1'h0};
  assign T_3418 = T_2933 ? tgts_T_3294_data : {{11'd0}, 1'h0};
  assign T_3420 = T_2934 ? tgts_T_3296_data : {{11'd0}, 1'h0};
  assign T_3422 = T_2935 ? tgts_T_3298_data : {{11'd0}, 1'h0};
  assign T_3424 = T_2936 ? tgts_T_3300_data : {{11'd0}, 1'h0};
  assign T_3426 = T_2937 ? tgts_T_3302_data : {{11'd0}, 1'h0};
  assign T_3428 = T_2938 ? tgts_T_3304_data : {{11'd0}, 1'h0};
  assign T_3430 = T_2939 ? tgts_T_3306_data : {{11'd0}, 1'h0};
  assign T_3432 = T_2940 ? tgts_T_3308_data : {{11'd0}, 1'h0};
  assign T_3434 = T_2941 ? tgts_T_3310_data : {{11'd0}, 1'h0};
  assign T_3436 = T_2942 ? tgts_T_3312_data : {{11'd0}, 1'h0};
  assign T_3438 = T_2943 ? tgts_T_3314_data : {{11'd0}, 1'h0};
  assign T_3440 = T_2944 ? tgts_T_3316_data : {{11'd0}, 1'h0};
  assign T_3442 = T_2945 ? tgts_T_3318_data : {{11'd0}, 1'h0};
  assign T_3444 = T_2946 ? tgts_T_3320_data : {{11'd0}, 1'h0};
  assign T_3446 = T_2947 ? tgts_T_3322_data : {{11'd0}, 1'h0};
  assign T_3448 = T_2948 ? tgts_T_3324_data : {{11'd0}, 1'h0};
  assign T_3450 = T_2949 ? tgts_T_3326_data : {{11'd0}, 1'h0};
  assign T_3452 = T_2950 ? tgts_T_3328_data : {{11'd0}, 1'h0};
  assign T_3454 = T_2951 ? tgts_T_3330_data : {{11'd0}, 1'h0};
  assign T_3456 = T_2952 ? tgts_T_3332_data : {{11'd0}, 1'h0};
  assign T_3458 = T_2953 ? tgts_T_3334_data : {{11'd0}, 1'h0};
  assign T_3460 = T_2954 ? tgts_T_3336_data : {{11'd0}, 1'h0};
  assign T_3462 = T_2955 ? tgts_T_3338_data : {{11'd0}, 1'h0};
  assign T_3464 = T_2956 ? tgts_T_3340_data : {{11'd0}, 1'h0};
  assign T_3466 = T_2957 ? tgts_T_3342_data : {{11'd0}, 1'h0};
  assign T_3468 = T_2958 ? tgts_T_3344_data : {{11'd0}, 1'h0};
  assign T_3470 = T_2959 ? tgts_T_3346_data : {{11'd0}, 1'h0};
  assign T_3472 = T_2960 ? tgts_T_3348_data : {{11'd0}, 1'h0};
  assign T_3474 = T_2961 ? tgts_T_3350_data : {{11'd0}, 1'h0};
  assign T_3476 = T_2962 ? tgts_T_3352_data : {{11'd0}, 1'h0};
  assign T_3478 = T_2963 ? tgts_T_3354_data : {{11'd0}, 1'h0};
  assign T_3480 = T_2964 ? tgts_T_3356_data : {{11'd0}, 1'h0};
  assign T_3482 = T_2965 ? tgts_T_3358_data : {{11'd0}, 1'h0};
  assign T_3484 = T_2966 ? tgts_T_3360_data : {{11'd0}, 1'h0};
  assign T_3486 = T_2967 ? tgts_T_3362_data : {{11'd0}, 1'h0};
  assign T_3488 = T_2968 ? tgts_T_3364_data : {{11'd0}, 1'h0};
  assign T_3490 = T_2969 ? tgts_T_3366_data : {{11'd0}, 1'h0};
  assign T_3492 = T_2970 ? tgts_T_3368_data : {{11'd0}, 1'h0};
  assign T_3494 = T_2971 ? tgts_T_3370_data : {{11'd0}, 1'h0};
  assign T_3496 = T_2972 ? tgts_T_3372_data : {{11'd0}, 1'h0};
  assign T_3498 = T_2973 ? tgts_T_3374_data : {{11'd0}, 1'h0};
  assign T_3500 = T_2974 ? tgts_T_3376_data : {{11'd0}, 1'h0};
  assign T_3502 = T_2975 ? tgts_T_3378_data : {{11'd0}, 1'h0};
  assign T_3504 = T_2976 ? tgts_T_3380_data : {{11'd0}, 1'h0};
  assign T_3506 = T_2977 ? tgts_T_3382_data : {{11'd0}, 1'h0};
  assign T_3508 = T_2978 ? tgts_T_3384_data : {{11'd0}, 1'h0};
  assign T_3510 = T_2979 ? tgts_T_3386_data : {{11'd0}, 1'h0};
  assign T_3512 = T_2980 ? tgts_T_3388_data : {{11'd0}, 1'h0};
  assign T_3514 = T_2981 ? tgts_T_3390_data : {{11'd0}, 1'h0};
  assign T_3516 = T_2982 ? tgts_T_3392_data : {{11'd0}, 1'h0};
  assign T_3518 = T_3394 | T_3396;
  assign T_3519 = T_3518 | T_3398;
  assign T_3520 = T_3519 | T_3400;
  assign T_3521 = T_3520 | T_3402;
  assign T_3522 = T_3521 | T_3404;
  assign T_3523 = T_3522 | T_3406;
  assign T_3524 = T_3523 | T_3408;
  assign T_3525 = T_3524 | T_3410;
  assign T_3526 = T_3525 | T_3412;
  assign T_3527 = T_3526 | T_3414;
  assign T_3528 = T_3527 | T_3416;
  assign T_3529 = T_3528 | T_3418;
  assign T_3530 = T_3529 | T_3420;
  assign T_3531 = T_3530 | T_3422;
  assign T_3532 = T_3531 | T_3424;
  assign T_3533 = T_3532 | T_3426;
  assign T_3534 = T_3533 | T_3428;
  assign T_3535 = T_3534 | T_3430;
  assign T_3536 = T_3535 | T_3432;
  assign T_3537 = T_3536 | T_3434;
  assign T_3538 = T_3537 | T_3436;
  assign T_3539 = T_3538 | T_3438;
  assign T_3540 = T_3539 | T_3440;
  assign T_3541 = T_3540 | T_3442;
  assign T_3542 = T_3541 | T_3444;
  assign T_3543 = T_3542 | T_3446;
  assign T_3544 = T_3543 | T_3448;
  assign T_3545 = T_3544 | T_3450;
  assign T_3546 = T_3545 | T_3452;
  assign T_3547 = T_3546 | T_3454;
  assign T_3548 = T_3547 | T_3456;
  assign T_3549 = T_3548 | T_3458;
  assign T_3550 = T_3549 | T_3460;
  assign T_3551 = T_3550 | T_3462;
  assign T_3552 = T_3551 | T_3464;
  assign T_3553 = T_3552 | T_3466;
  assign T_3554 = T_3553 | T_3468;
  assign T_3555 = T_3554 | T_3470;
  assign T_3556 = T_3555 | T_3472;
  assign T_3557 = T_3556 | T_3474;
  assign T_3558 = T_3557 | T_3476;
  assign T_3559 = T_3558 | T_3478;
  assign T_3560 = T_3559 | T_3480;
  assign T_3561 = T_3560 | T_3482;
  assign T_3562 = T_3561 | T_3484;
  assign T_3563 = T_3562 | T_3486;
  assign T_3564 = T_3563 | T_3488;
  assign T_3565 = T_3564 | T_3490;
  assign T_3566 = T_3565 | T_3492;
  assign T_3567 = T_3566 | T_3494;
  assign T_3568 = T_3567 | T_3496;
  assign T_3569 = T_3568 | T_3498;
  assign T_3570 = T_3569 | T_3500;
  assign T_3571 = T_3570 | T_3502;
  assign T_3572 = T_3571 | T_3504;
  assign T_3573 = T_3572 | T_3506;
  assign T_3574 = T_3573 | T_3508;
  assign T_3575 = T_3574 | T_3510;
  assign T_3576 = T_3575 | T_3512;
  assign T_3577 = T_3576 | T_3514;
  assign T_3578 = T_3577 | T_3516;
  assign T_3579 = T_3578;
  assign T_3580 = {T_3206,T_3579};
  assign T_3581 = hits[61:32];
  assign T_3582 = hits[31:0];
  assign GEN_848 = {{29'd0}, 1'h0};
  assign T_3584 = T_3581 != GEN_848;
  assign GEN_849 = {{2'd0}, T_3581};
  assign T_3585 = GEN_849 | T_3582;
  assign T_3586 = T_3585[31:16];
  assign T_3587 = T_3585[15:0];
  assign GEN_850 = {{15'd0}, 1'h0};
  assign T_3589 = T_3586 != GEN_850;
  assign T_3590 = T_3586 | T_3587;
  assign T_3591 = T_3590[15:8];
  assign T_3592 = T_3590[7:0];
  assign GEN_851 = {{7'd0}, 1'h0};
  assign T_3594 = T_3591 != GEN_851;
  assign T_3595 = T_3591 | T_3592;
  assign T_3596 = T_3595[7:4];
  assign T_3597 = T_3595[3:0];
  assign GEN_852 = {{3'd0}, 1'h0};
  assign T_3599 = T_3596 != GEN_852;
  assign T_3600 = T_3596 | T_3597;
  assign T_3601 = T_3600[3:2];
  assign T_3602 = T_3600[1:0];
  assign T_3604 = T_3601 != GEN_707;
  assign T_3605 = T_3601 | T_3602;
  assign T_3606 = T_3605[1];
  assign T_3607 = {T_3604,T_3606};
  assign T_3608 = {T_3599,T_3607};
  assign T_3609 = {T_3594,T_3608};
  assign T_3610 = {T_3589,T_3609};
  assign T_3611 = {T_3584,T_3610};
  assign T_3616_T_3942_addr = T_3941;
  assign T_3616_T_3942_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_3616_T_3942_data = T_3616[T_3616_T_3942_addr];
  `else
  assign T_3616_T_3942_data = T_3616_T_3942_addr >= 8'h80 ? $random : T_3616[T_3616_T_3942_addr];
  `endif
  assign T_3616_T_3949_data = T_3958;
  assign T_3616_T_3949_addr = T_3948;
  assign T_3616_T_3949_mask = T_3946;
  assign T_3616_T_3949_en = T_3946;
  assign T_3683 = T_2921 ? isJump_0 : 1'h0;
  assign T_3686 = T_2922 ? isJump_1 : 1'h0;
  assign T_3689 = T_2923 ? isJump_2 : 1'h0;
  assign T_3692 = T_2924 ? isJump_3 : 1'h0;
  assign T_3695 = T_2925 ? isJump_4 : 1'h0;
  assign T_3698 = T_2926 ? isJump_5 : 1'h0;
  assign T_3701 = T_2927 ? isJump_6 : 1'h0;
  assign T_3704 = T_2928 ? isJump_7 : 1'h0;
  assign T_3707 = T_2929 ? isJump_8 : 1'h0;
  assign T_3710 = T_2930 ? isJump_9 : 1'h0;
  assign T_3713 = T_2931 ? isJump_10 : 1'h0;
  assign T_3716 = T_2932 ? isJump_11 : 1'h0;
  assign T_3719 = T_2933 ? isJump_12 : 1'h0;
  assign T_3722 = T_2934 ? isJump_13 : 1'h0;
  assign T_3725 = T_2935 ? isJump_14 : 1'h0;
  assign T_3728 = T_2936 ? isJump_15 : 1'h0;
  assign T_3731 = T_2937 ? isJump_16 : 1'h0;
  assign T_3734 = T_2938 ? isJump_17 : 1'h0;
  assign T_3737 = T_2939 ? isJump_18 : 1'h0;
  assign T_3740 = T_2940 ? isJump_19 : 1'h0;
  assign T_3743 = T_2941 ? isJump_20 : 1'h0;
  assign T_3746 = T_2942 ? isJump_21 : 1'h0;
  assign T_3749 = T_2943 ? isJump_22 : 1'h0;
  assign T_3752 = T_2944 ? isJump_23 : 1'h0;
  assign T_3755 = T_2945 ? isJump_24 : 1'h0;
  assign T_3758 = T_2946 ? isJump_25 : 1'h0;
  assign T_3761 = T_2947 ? isJump_26 : 1'h0;
  assign T_3764 = T_2948 ? isJump_27 : 1'h0;
  assign T_3767 = T_2949 ? isJump_28 : 1'h0;
  assign T_3770 = T_2950 ? isJump_29 : 1'h0;
  assign T_3773 = T_2951 ? isJump_30 : 1'h0;
  assign T_3776 = T_2952 ? isJump_31 : 1'h0;
  assign T_3779 = T_2953 ? isJump_32 : 1'h0;
  assign T_3782 = T_2954 ? isJump_33 : 1'h0;
  assign T_3785 = T_2955 ? isJump_34 : 1'h0;
  assign T_3788 = T_2956 ? isJump_35 : 1'h0;
  assign T_3791 = T_2957 ? isJump_36 : 1'h0;
  assign T_3794 = T_2958 ? isJump_37 : 1'h0;
  assign T_3797 = T_2959 ? isJump_38 : 1'h0;
  assign T_3800 = T_2960 ? isJump_39 : 1'h0;
  assign T_3803 = T_2961 ? isJump_40 : 1'h0;
  assign T_3806 = T_2962 ? isJump_41 : 1'h0;
  assign T_3809 = T_2963 ? isJump_42 : 1'h0;
  assign T_3812 = T_2964 ? isJump_43 : 1'h0;
  assign T_3815 = T_2965 ? isJump_44 : 1'h0;
  assign T_3818 = T_2966 ? isJump_45 : 1'h0;
  assign T_3821 = T_2967 ? isJump_46 : 1'h0;
  assign T_3824 = T_2968 ? isJump_47 : 1'h0;
  assign T_3827 = T_2969 ? isJump_48 : 1'h0;
  assign T_3830 = T_2970 ? isJump_49 : 1'h0;
  assign T_3833 = T_2971 ? isJump_50 : 1'h0;
  assign T_3836 = T_2972 ? isJump_51 : 1'h0;
  assign T_3839 = T_2973 ? isJump_52 : 1'h0;
  assign T_3842 = T_2974 ? isJump_53 : 1'h0;
  assign T_3845 = T_2975 ? isJump_54 : 1'h0;
  assign T_3848 = T_2976 ? isJump_55 : 1'h0;
  assign T_3851 = T_2977 ? isJump_56 : 1'h0;
  assign T_3854 = T_2978 ? isJump_57 : 1'h0;
  assign T_3857 = T_2979 ? isJump_58 : 1'h0;
  assign T_3860 = T_2980 ? isJump_59 : 1'h0;
  assign T_3863 = T_2981 ? isJump_60 : 1'h0;
  assign T_3866 = T_2982 ? isJump_61 : 1'h0;
  assign T_3868 = T_3683 | T_3686;
  assign T_3869 = T_3868 | T_3689;
  assign T_3870 = T_3869 | T_3692;
  assign T_3871 = T_3870 | T_3695;
  assign T_3872 = T_3871 | T_3698;
  assign T_3873 = T_3872 | T_3701;
  assign T_3874 = T_3873 | T_3704;
  assign T_3875 = T_3874 | T_3707;
  assign T_3876 = T_3875 | T_3710;
  assign T_3877 = T_3876 | T_3713;
  assign T_3878 = T_3877 | T_3716;
  assign T_3879 = T_3878 | T_3719;
  assign T_3880 = T_3879 | T_3722;
  assign T_3881 = T_3880 | T_3725;
  assign T_3882 = T_3881 | T_3728;
  assign T_3883 = T_3882 | T_3731;
  assign T_3884 = T_3883 | T_3734;
  assign T_3885 = T_3884 | T_3737;
  assign T_3886 = T_3885 | T_3740;
  assign T_3887 = T_3886 | T_3743;
  assign T_3888 = T_3887 | T_3746;
  assign T_3889 = T_3888 | T_3749;
  assign T_3890 = T_3889 | T_3752;
  assign T_3891 = T_3890 | T_3755;
  assign T_3892 = T_3891 | T_3758;
  assign T_3893 = T_3892 | T_3761;
  assign T_3894 = T_3893 | T_3764;
  assign T_3895 = T_3894 | T_3767;
  assign T_3896 = T_3895 | T_3770;
  assign T_3897 = T_3896 | T_3773;
  assign T_3898 = T_3897 | T_3776;
  assign T_3899 = T_3898 | T_3779;
  assign T_3900 = T_3899 | T_3782;
  assign T_3901 = T_3900 | T_3785;
  assign T_3902 = T_3901 | T_3788;
  assign T_3903 = T_3902 | T_3791;
  assign T_3904 = T_3903 | T_3794;
  assign T_3905 = T_3904 | T_3797;
  assign T_3906 = T_3905 | T_3800;
  assign T_3907 = T_3906 | T_3803;
  assign T_3908 = T_3907 | T_3806;
  assign T_3909 = T_3908 | T_3809;
  assign T_3910 = T_3909 | T_3812;
  assign T_3911 = T_3910 | T_3815;
  assign T_3912 = T_3911 | T_3818;
  assign T_3913 = T_3912 | T_3821;
  assign T_3914 = T_3913 | T_3824;
  assign T_3915 = T_3914 | T_3827;
  assign T_3916 = T_3915 | T_3830;
  assign T_3917 = T_3916 | T_3833;
  assign T_3918 = T_3917 | T_3836;
  assign T_3919 = T_3918 | T_3839;
  assign T_3920 = T_3919 | T_3842;
  assign T_3921 = T_3920 | T_3845;
  assign T_3922 = T_3921 | T_3848;
  assign T_3923 = T_3922 | T_3851;
  assign T_3924 = T_3923 | T_3854;
  assign T_3925 = T_3924 | T_3857;
  assign T_3926 = T_3925 | T_3860;
  assign T_3927 = T_3926 | T_3863;
  assign T_3928 = T_3927 | T_3866;
  assign T_3929 = T_3928;
  assign T_3931 = T_3929 == 1'h0;
  assign T_3932 = io_req_valid & io_resp_valid;
  assign T_3933 = T_3932 & T_3931;
  assign T_3937_history = T_3618;
  assign T_3937_value = T_3616_T_3942_data;
  assign T_3940 = io_req_bits_addr[8:2];
  assign T_3941 = T_3940 ^ T_3618;
  assign T_3943 = T_3937_value[0];
  assign T_3944 = T_3618[6:1];
  assign T_3945 = {T_3943,T_3944};
  assign GEN_424 = T_3933 ? T_3945 : T_3618;
  assign T_3946 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T_3947 = io_bht_update_bits_pc[8:2];
  assign T_3948 = T_3947 ^ io_bht_update_bits_prediction_bits_bht_history;
  assign T_3950 = io_bht_update_bits_prediction_bits_bht_value[1];
  assign T_3951 = io_bht_update_bits_prediction_bits_bht_value[0];
  assign T_3952 = T_3950 & T_3951;
  assign T_3955 = T_3950 | T_3951;
  assign T_3956 = T_3955 & io_bht_update_bits_taken;
  assign T_3957 = T_3952 | T_3956;
  assign T_3958 = {io_bht_update_bits_taken,T_3957};
  assign T_3959 = io_bht_update_bits_prediction_bits_bht_history[6:1];
  assign T_3960 = {io_bht_update_bits_taken,T_3959};
  assign GEN_425 = io_bht_update_bits_mispredict ? T_3960 : GEN_424;
  assign GEN_431 = T_3946 ? GEN_425 : GEN_424;
  assign T_3963 = T_3943 == 1'h0;
  assign T_3964 = T_3963 & T_3931;
  assign GEN_432 = T_3964 ? 1'h0 : io_resp_valid;
  assign T_4042 = T_2921 ? useRAS_0 : 1'h0;
  assign T_4045 = T_2922 ? useRAS_1 : 1'h0;
  assign T_4048 = T_2923 ? useRAS_2 : 1'h0;
  assign T_4051 = T_2924 ? useRAS_3 : 1'h0;
  assign T_4054 = T_2925 ? useRAS_4 : 1'h0;
  assign T_4057 = T_2926 ? useRAS_5 : 1'h0;
  assign T_4060 = T_2927 ? useRAS_6 : 1'h0;
  assign T_4063 = T_2928 ? useRAS_7 : 1'h0;
  assign T_4066 = T_2929 ? useRAS_8 : 1'h0;
  assign T_4069 = T_2930 ? useRAS_9 : 1'h0;
  assign T_4072 = T_2931 ? useRAS_10 : 1'h0;
  assign T_4075 = T_2932 ? useRAS_11 : 1'h0;
  assign T_4078 = T_2933 ? useRAS_12 : 1'h0;
  assign T_4081 = T_2934 ? useRAS_13 : 1'h0;
  assign T_4084 = T_2935 ? useRAS_14 : 1'h0;
  assign T_4087 = T_2936 ? useRAS_15 : 1'h0;
  assign T_4090 = T_2937 ? useRAS_16 : 1'h0;
  assign T_4093 = T_2938 ? useRAS_17 : 1'h0;
  assign T_4096 = T_2939 ? useRAS_18 : 1'h0;
  assign T_4099 = T_2940 ? useRAS_19 : 1'h0;
  assign T_4102 = T_2941 ? useRAS_20 : 1'h0;
  assign T_4105 = T_2942 ? useRAS_21 : 1'h0;
  assign T_4108 = T_2943 ? useRAS_22 : 1'h0;
  assign T_4111 = T_2944 ? useRAS_23 : 1'h0;
  assign T_4114 = T_2945 ? useRAS_24 : 1'h0;
  assign T_4117 = T_2946 ? useRAS_25 : 1'h0;
  assign T_4120 = T_2947 ? useRAS_26 : 1'h0;
  assign T_4123 = T_2948 ? useRAS_27 : 1'h0;
  assign T_4126 = T_2949 ? useRAS_28 : 1'h0;
  assign T_4129 = T_2950 ? useRAS_29 : 1'h0;
  assign T_4132 = T_2951 ? useRAS_30 : 1'h0;
  assign T_4135 = T_2952 ? useRAS_31 : 1'h0;
  assign T_4138 = T_2953 ? useRAS_32 : 1'h0;
  assign T_4141 = T_2954 ? useRAS_33 : 1'h0;
  assign T_4144 = T_2955 ? useRAS_34 : 1'h0;
  assign T_4147 = T_2956 ? useRAS_35 : 1'h0;
  assign T_4150 = T_2957 ? useRAS_36 : 1'h0;
  assign T_4153 = T_2958 ? useRAS_37 : 1'h0;
  assign T_4156 = T_2959 ? useRAS_38 : 1'h0;
  assign T_4159 = T_2960 ? useRAS_39 : 1'h0;
  assign T_4162 = T_2961 ? useRAS_40 : 1'h0;
  assign T_4165 = T_2962 ? useRAS_41 : 1'h0;
  assign T_4168 = T_2963 ? useRAS_42 : 1'h0;
  assign T_4171 = T_2964 ? useRAS_43 : 1'h0;
  assign T_4174 = T_2965 ? useRAS_44 : 1'h0;
  assign T_4177 = T_2966 ? useRAS_45 : 1'h0;
  assign T_4180 = T_2967 ? useRAS_46 : 1'h0;
  assign T_4183 = T_2968 ? useRAS_47 : 1'h0;
  assign T_4186 = T_2969 ? useRAS_48 : 1'h0;
  assign T_4189 = T_2970 ? useRAS_49 : 1'h0;
  assign T_4192 = T_2971 ? useRAS_50 : 1'h0;
  assign T_4195 = T_2972 ? useRAS_51 : 1'h0;
  assign T_4198 = T_2973 ? useRAS_52 : 1'h0;
  assign T_4201 = T_2974 ? useRAS_53 : 1'h0;
  assign T_4204 = T_2975 ? useRAS_54 : 1'h0;
  assign T_4207 = T_2976 ? useRAS_55 : 1'h0;
  assign T_4210 = T_2977 ? useRAS_56 : 1'h0;
  assign T_4213 = T_2978 ? useRAS_57 : 1'h0;
  assign T_4216 = T_2979 ? useRAS_58 : 1'h0;
  assign T_4219 = T_2980 ? useRAS_59 : 1'h0;
  assign T_4222 = T_2981 ? useRAS_60 : 1'h0;
  assign T_4225 = T_2982 ? useRAS_61 : 1'h0;
  assign T_4227 = T_4042 | T_4045;
  assign T_4228 = T_4227 | T_4048;
  assign T_4229 = T_4228 | T_4051;
  assign T_4230 = T_4229 | T_4054;
  assign T_4231 = T_4230 | T_4057;
  assign T_4232 = T_4231 | T_4060;
  assign T_4233 = T_4232 | T_4063;
  assign T_4234 = T_4233 | T_4066;
  assign T_4235 = T_4234 | T_4069;
  assign T_4236 = T_4235 | T_4072;
  assign T_4237 = T_4236 | T_4075;
  assign T_4238 = T_4237 | T_4078;
  assign T_4239 = T_4238 | T_4081;
  assign T_4240 = T_4239 | T_4084;
  assign T_4241 = T_4240 | T_4087;
  assign T_4242 = T_4241 | T_4090;
  assign T_4243 = T_4242 | T_4093;
  assign T_4244 = T_4243 | T_4096;
  assign T_4245 = T_4244 | T_4099;
  assign T_4246 = T_4245 | T_4102;
  assign T_4247 = T_4246 | T_4105;
  assign T_4248 = T_4247 | T_4108;
  assign T_4249 = T_4248 | T_4111;
  assign T_4250 = T_4249 | T_4114;
  assign T_4251 = T_4250 | T_4117;
  assign T_4252 = T_4251 | T_4120;
  assign T_4253 = T_4252 | T_4123;
  assign T_4254 = T_4253 | T_4126;
  assign T_4255 = T_4254 | T_4129;
  assign T_4256 = T_4255 | T_4132;
  assign T_4257 = T_4256 | T_4135;
  assign T_4258 = T_4257 | T_4138;
  assign T_4259 = T_4258 | T_4141;
  assign T_4260 = T_4259 | T_4144;
  assign T_4261 = T_4260 | T_4147;
  assign T_4262 = T_4261 | T_4150;
  assign T_4263 = T_4262 | T_4153;
  assign T_4264 = T_4263 | T_4156;
  assign T_4265 = T_4264 | T_4159;
  assign T_4266 = T_4265 | T_4162;
  assign T_4267 = T_4266 | T_4165;
  assign T_4268 = T_4267 | T_4168;
  assign T_4269 = T_4268 | T_4171;
  assign T_4270 = T_4269 | T_4174;
  assign T_4271 = T_4270 | T_4177;
  assign T_4272 = T_4271 | T_4180;
  assign T_4273 = T_4272 | T_4183;
  assign T_4274 = T_4273 | T_4186;
  assign T_4275 = T_4274 | T_4189;
  assign T_4276 = T_4275 | T_4192;
  assign T_4277 = T_4276 | T_4195;
  assign T_4278 = T_4277 | T_4198;
  assign T_4279 = T_4278 | T_4201;
  assign T_4280 = T_4279 | T_4204;
  assign T_4281 = T_4280 | T_4207;
  assign T_4282 = T_4281 | T_4210;
  assign T_4283 = T_4282 | T_4213;
  assign T_4284 = T_4283 | T_4216;
  assign T_4285 = T_4284 | T_4219;
  assign T_4286 = T_4285 | T_4222;
  assign T_4287 = T_4286 | T_4225;
  assign T_4288 = T_4287;
  assign T_4290 = T_3967 == GEN_707;
  assign T_4292 = T_4290 == 1'h0;
  assign T_4293 = T_4292 & T_4288;
  assign GEN_2 = GEN_433;
  assign GEN_433 = T_3969 ? T_3976_1 : T_3976_0;
  assign GEN_435 = T_4293 ? GEN_2 : T_3580;
  assign T_4295 = T_3967 < 2'h2;
  assign GEN_855 = {{1'd0}, 1'h1};
  assign T_4297 = T_3967 + GEN_855;
  assign T_4298 = T_4297[1:0];
  assign GEN_436 = T_4295 ? T_4298 : T_3967;
  assign T_4304 = T_3969 + 1'h1;
  assign T_4305 = T_4304[0:0];
  assign GEN_3 = io_ras_update_bits_returnAddr;
  assign GEN_437 = 1'h0 == T_4305 ? GEN_3 : T_3976_0;
  assign GEN_438 = T_4305 ? GEN_3 : T_3976_1;
  assign GEN_439 = T_4288 ? io_ras_update_bits_returnAddr : GEN_435;
  assign GEN_440 = io_ras_update_bits_isCall ? GEN_436 : T_3967;
  assign GEN_442 = io_ras_update_bits_isCall ? GEN_437 : T_3976_0;
  assign GEN_443 = io_ras_update_bits_isCall ? GEN_438 : T_3976_1;
  assign GEN_444 = io_ras_update_bits_isCall ? T_4305 : T_3969;
  assign GEN_445 = io_ras_update_bits_isCall ? GEN_439 : GEN_435;
  assign T_4308 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T_4310 = io_ras_update_bits_isCall == 1'h0;
  assign T_4311 = T_4310 & T_4308;
  assign T_4317 = T_3967 - GEN_855;
  assign T_4318 = T_4317[1:0];
  assign T_4324 = T_3969 - 1'h1;
  assign T_4325 = T_4324[0:0];
  assign GEN_446 = T_4292 ? T_4318 : GEN_440;
  assign GEN_447 = T_4292 ? T_4325 : GEN_444;
  assign GEN_448 = T_4311 ? GEN_446 : GEN_440;
  assign GEN_449 = T_4311 ? GEN_447 : GEN_444;
  assign GEN_450 = io_ras_update_valid ? GEN_448 : T_3967;
  assign GEN_452 = io_ras_update_valid ? GEN_442 : T_3976_0;
  assign GEN_453 = io_ras_update_valid ? GEN_443 : T_3976_1;
  assign GEN_454 = io_ras_update_valid ? GEN_449 : T_3969;
  assign GEN_455 = io_ras_update_valid ? GEN_445 : GEN_435;
  assign GEN_456 = io_invalidate ? {{1'd0}, 1'h0} : GEN_450;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_146 = {2{$random}};
  idxValid = GEN_146[61:0];
  GEN_147 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    idxs[initvar] = GEN_147[11:0];
  GEN_148 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    idxPages[initvar] = GEN_148[2:0];
  GEN_149 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    tgts[initvar] = GEN_149[11:0];
  GEN_150 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    tgtPages[initvar] = GEN_150[2:0];
  GEN_151 = {1{$random}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    pages[initvar] = GEN_151[26:0];
  GEN_152 = {1{$random}};
  pageValid = GEN_152[5:0];
  GEN_153 = {1{$random}};
  useRAS_0 = GEN_153[0:0];
  GEN_154 = {1{$random}};
  useRAS_1 = GEN_154[0:0];
  GEN_155 = {1{$random}};
  useRAS_2 = GEN_155[0:0];
  GEN_156 = {1{$random}};
  useRAS_3 = GEN_156[0:0];
  GEN_157 = {1{$random}};
  useRAS_4 = GEN_157[0:0];
  GEN_158 = {1{$random}};
  useRAS_5 = GEN_158[0:0];
  GEN_159 = {1{$random}};
  useRAS_6 = GEN_159[0:0];
  GEN_160 = {1{$random}};
  useRAS_7 = GEN_160[0:0];
  GEN_161 = {1{$random}};
  useRAS_8 = GEN_161[0:0];
  GEN_162 = {1{$random}};
  useRAS_9 = GEN_162[0:0];
  GEN_163 = {1{$random}};
  useRAS_10 = GEN_163[0:0];
  GEN_164 = {1{$random}};
  useRAS_11 = GEN_164[0:0];
  GEN_165 = {1{$random}};
  useRAS_12 = GEN_165[0:0];
  GEN_166 = {1{$random}};
  useRAS_13 = GEN_166[0:0];
  GEN_167 = {1{$random}};
  useRAS_14 = GEN_167[0:0];
  GEN_168 = {1{$random}};
  useRAS_15 = GEN_168[0:0];
  GEN_169 = {1{$random}};
  useRAS_16 = GEN_169[0:0];
  GEN_170 = {1{$random}};
  useRAS_17 = GEN_170[0:0];
  GEN_171 = {1{$random}};
  useRAS_18 = GEN_171[0:0];
  GEN_172 = {1{$random}};
  useRAS_19 = GEN_172[0:0];
  GEN_173 = {1{$random}};
  useRAS_20 = GEN_173[0:0];
  GEN_174 = {1{$random}};
  useRAS_21 = GEN_174[0:0];
  GEN_175 = {1{$random}};
  useRAS_22 = GEN_175[0:0];
  GEN_177 = {1{$random}};
  useRAS_23 = GEN_177[0:0];
  GEN_178 = {1{$random}};
  useRAS_24 = GEN_178[0:0];
  GEN_179 = {1{$random}};
  useRAS_25 = GEN_179[0:0];
  GEN_180 = {1{$random}};
  useRAS_26 = GEN_180[0:0];
  GEN_181 = {1{$random}};
  useRAS_27 = GEN_181[0:0];
  GEN_182 = {1{$random}};
  useRAS_28 = GEN_182[0:0];
  GEN_183 = {1{$random}};
  useRAS_29 = GEN_183[0:0];
  GEN_184 = {1{$random}};
  useRAS_30 = GEN_184[0:0];
  GEN_185 = {1{$random}};
  useRAS_31 = GEN_185[0:0];
  GEN_186 = {1{$random}};
  useRAS_32 = GEN_186[0:0];
  GEN_187 = {1{$random}};
  useRAS_33 = GEN_187[0:0];
  GEN_188 = {1{$random}};
  useRAS_34 = GEN_188[0:0];
  GEN_189 = {1{$random}};
  useRAS_35 = GEN_189[0:0];
  GEN_190 = {1{$random}};
  useRAS_36 = GEN_190[0:0];
  GEN_191 = {1{$random}};
  useRAS_37 = GEN_191[0:0];
  GEN_192 = {1{$random}};
  useRAS_38 = GEN_192[0:0];
  GEN_193 = {1{$random}};
  useRAS_39 = GEN_193[0:0];
  GEN_194 = {1{$random}};
  useRAS_40 = GEN_194[0:0];
  GEN_195 = {1{$random}};
  useRAS_41 = GEN_195[0:0];
  GEN_196 = {1{$random}};
  useRAS_42 = GEN_196[0:0];
  GEN_197 = {1{$random}};
  useRAS_43 = GEN_197[0:0];
  GEN_198 = {1{$random}};
  useRAS_44 = GEN_198[0:0];
  GEN_199 = {1{$random}};
  useRAS_45 = GEN_199[0:0];
  GEN_200 = {1{$random}};
  useRAS_46 = GEN_200[0:0];
  GEN_201 = {1{$random}};
  useRAS_47 = GEN_201[0:0];
  GEN_202 = {1{$random}};
  useRAS_48 = GEN_202[0:0];
  GEN_203 = {1{$random}};
  useRAS_49 = GEN_203[0:0];
  GEN_204 = {1{$random}};
  useRAS_50 = GEN_204[0:0];
  GEN_205 = {1{$random}};
  useRAS_51 = GEN_205[0:0];
  GEN_206 = {1{$random}};
  useRAS_52 = GEN_206[0:0];
  GEN_207 = {1{$random}};
  useRAS_53 = GEN_207[0:0];
  GEN_208 = {1{$random}};
  useRAS_54 = GEN_208[0:0];
  GEN_209 = {1{$random}};
  useRAS_55 = GEN_209[0:0];
  GEN_210 = {1{$random}};
  useRAS_56 = GEN_210[0:0];
  GEN_211 = {1{$random}};
  useRAS_57 = GEN_211[0:0];
  GEN_212 = {1{$random}};
  useRAS_58 = GEN_212[0:0];
  GEN_213 = {1{$random}};
  useRAS_59 = GEN_213[0:0];
  GEN_214 = {1{$random}};
  useRAS_60 = GEN_214[0:0];
  GEN_215 = {1{$random}};
  useRAS_61 = GEN_215[0:0];
  GEN_216 = {1{$random}};
  isJump_0 = GEN_216[0:0];
  GEN_217 = {1{$random}};
  isJump_1 = GEN_217[0:0];
  GEN_218 = {1{$random}};
  isJump_2 = GEN_218[0:0];
  GEN_219 = {1{$random}};
  isJump_3 = GEN_219[0:0];
  GEN_220 = {1{$random}};
  isJump_4 = GEN_220[0:0];
  GEN_221 = {1{$random}};
  isJump_5 = GEN_221[0:0];
  GEN_222 = {1{$random}};
  isJump_6 = GEN_222[0:0];
  GEN_223 = {1{$random}};
  isJump_7 = GEN_223[0:0];
  GEN_224 = {1{$random}};
  isJump_8 = GEN_224[0:0];
  GEN_225 = {1{$random}};
  isJump_9 = GEN_225[0:0];
  GEN_226 = {1{$random}};
  isJump_10 = GEN_226[0:0];
  GEN_227 = {1{$random}};
  isJump_11 = GEN_227[0:0];
  GEN_228 = {1{$random}};
  isJump_12 = GEN_228[0:0];
  GEN_229 = {1{$random}};
  isJump_13 = GEN_229[0:0];
  GEN_230 = {1{$random}};
  isJump_14 = GEN_230[0:0];
  GEN_231 = {1{$random}};
  isJump_15 = GEN_231[0:0];
  GEN_232 = {1{$random}};
  isJump_16 = GEN_232[0:0];
  GEN_233 = {1{$random}};
  isJump_17 = GEN_233[0:0];
  GEN_234 = {1{$random}};
  isJump_18 = GEN_234[0:0];
  GEN_235 = {1{$random}};
  isJump_19 = GEN_235[0:0];
  GEN_236 = {1{$random}};
  isJump_20 = GEN_236[0:0];
  GEN_237 = {1{$random}};
  isJump_21 = GEN_237[0:0];
  GEN_238 = {1{$random}};
  isJump_22 = GEN_238[0:0];
  GEN_240 = {1{$random}};
  isJump_23 = GEN_240[0:0];
  GEN_241 = {1{$random}};
  isJump_24 = GEN_241[0:0];
  GEN_242 = {1{$random}};
  isJump_25 = GEN_242[0:0];
  GEN_243 = {1{$random}};
  isJump_26 = GEN_243[0:0];
  GEN_244 = {1{$random}};
  isJump_27 = GEN_244[0:0];
  GEN_245 = {1{$random}};
  isJump_28 = GEN_245[0:0];
  GEN_246 = {1{$random}};
  isJump_29 = GEN_246[0:0];
  GEN_247 = {1{$random}};
  isJump_30 = GEN_247[0:0];
  GEN_248 = {1{$random}};
  isJump_31 = GEN_248[0:0];
  GEN_249 = {1{$random}};
  isJump_32 = GEN_249[0:0];
  GEN_250 = {1{$random}};
  isJump_33 = GEN_250[0:0];
  GEN_251 = {1{$random}};
  isJump_34 = GEN_251[0:0];
  GEN_252 = {1{$random}};
  isJump_35 = GEN_252[0:0];
  GEN_253 = {1{$random}};
  isJump_36 = GEN_253[0:0];
  GEN_254 = {1{$random}};
  isJump_37 = GEN_254[0:0];
  GEN_255 = {1{$random}};
  isJump_38 = GEN_255[0:0];
  GEN_256 = {1{$random}};
  isJump_39 = GEN_256[0:0];
  GEN_257 = {1{$random}};
  isJump_40 = GEN_257[0:0];
  GEN_258 = {1{$random}};
  isJump_41 = GEN_258[0:0];
  GEN_259 = {1{$random}};
  isJump_42 = GEN_259[0:0];
  GEN_260 = {1{$random}};
  isJump_43 = GEN_260[0:0];
  GEN_323 = {1{$random}};
  isJump_44 = GEN_323[0:0];
  GEN_386 = {1{$random}};
  isJump_45 = GEN_386[0:0];
  GEN_387 = {1{$random}};
  isJump_46 = GEN_387[0:0];
  GEN_388 = {1{$random}};
  isJump_47 = GEN_388[0:0];
  GEN_389 = {1{$random}};
  isJump_48 = GEN_389[0:0];
  GEN_390 = {1{$random}};
  isJump_49 = GEN_390[0:0];
  GEN_391 = {1{$random}};
  isJump_50 = GEN_391[0:0];
  GEN_392 = {1{$random}};
  isJump_51 = GEN_392[0:0];
  GEN_394 = {1{$random}};
  isJump_52 = GEN_394[0:0];
  GEN_395 = {1{$random}};
  isJump_53 = GEN_395[0:0];
  GEN_396 = {1{$random}};
  isJump_54 = GEN_396[0:0];
  GEN_397 = {1{$random}};
  isJump_55 = GEN_397[0:0];
  GEN_399 = {1{$random}};
  isJump_56 = GEN_399[0:0];
  GEN_400 = {1{$random}};
  isJump_57 = GEN_400[0:0];
  GEN_401 = {1{$random}};
  isJump_58 = GEN_401[0:0];
  GEN_402 = {1{$random}};
  isJump_59 = GEN_402[0:0];
  GEN_404 = {1{$random}};
  isJump_60 = GEN_404[0:0];
  GEN_405 = {1{$random}};
  isJump_61 = GEN_405[0:0];
  GEN_406 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    brIdx[initvar] = GEN_406[0:0];
  GEN_407 = {1{$random}};
  T_1215 = GEN_407[0:0];
  GEN_409 = {1{$random}};
  T_1216_prediction_valid = GEN_409[0:0];
  GEN_410 = {1{$random}};
  T_1216_prediction_bits_taken = GEN_410[0:0];
  GEN_411 = {1{$random}};
  T_1216_prediction_bits_mask = GEN_411[0:0];
  GEN_412 = {1{$random}};
  T_1216_prediction_bits_bridx = GEN_412[0:0];
  GEN_414 = {2{$random}};
  T_1216_prediction_bits_target = GEN_414[38:0];
  GEN_415 = {1{$random}};
  T_1216_prediction_bits_entry = GEN_415[5:0];
  GEN_416 = {1{$random}};
  T_1216_prediction_bits_bht_history = GEN_416[6:0];
  GEN_417 = {1{$random}};
  T_1216_prediction_bits_bht_value = GEN_417[1:0];
  GEN_419 = {2{$random}};
  T_1216_pc = GEN_419[38:0];
  GEN_420 = {2{$random}};
  T_1216_target = GEN_420[38:0];
  GEN_426 = {1{$random}};
  T_1216_taken = GEN_426[0:0];
  GEN_427 = {1{$random}};
  T_1216_isJump = GEN_427[0:0];
  GEN_428 = {1{$random}};
  T_1216_isReturn = GEN_428[0:0];
  GEN_429 = {2{$random}};
  T_1216_br_pc = GEN_429[38:0];
  GEN_430 = {1{$random}};
  nextRepl = GEN_430[5:0];
  GEN_434 = {1{$random}};
  T_2536 = GEN_434[2:0];
  GEN_441 = {1{$random}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    T_3616[initvar] = GEN_441[1:0];
  GEN_451 = {1{$random}};
  T_3618 = GEN_451[6:0];
  GEN_458 = {1{$random}};
  T_3967 = GEN_458[1:0];
  GEN_459 = {1{$random}};
  T_3969 = GEN_459[0:0];
  GEN_460 = {2{$random}};
  T_3976_0 = GEN_460[38:0];
  GEN_461 = {2{$random}};
  T_3976_1 = GEN_461[38:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      idxValid <= 62'h0;
    end else begin
      idxValid <= GEN_422[61:0];
    end
    if(idxs_T_2872_en & idxs_T_2872_mask) begin
      idxs[idxs_T_2872_addr] <= idxs_T_2872_data;
    end
    if(idxPages_T_2874_en & idxPages_T_2874_mask) begin
      idxPages[idxPages_T_2874_addr] <= idxPages_T_2874_data;
    end
    if(tgts_T_2873_en & tgts_T_2873_mask) begin
      tgts[tgts_T_2873_addr] <= tgts_T_2873_data;
    end
    if(tgtPages_T_2875_en & tgtPages_T_2875_mask) begin
      tgtPages[tgtPages_T_2875_addr] <= tgtPages_T_2875_data;
    end
    if(pages_T_2891_en & pages_T_2891_mask) begin
      pages[pages_T_2891_addr] <= pages_T_2891_data;
    end
    if(pages_T_2895_en & pages_T_2895_mask) begin
      pages[pages_T_2895_addr] <= pages_T_2895_data;
    end
    if(pages_T_2899_en & pages_T_2899_mask) begin
      pages[pages_T_2899_addr] <= pages_T_2899_data;
    end
    if(pages_T_2907_en & pages_T_2907_mask) begin
      pages[pages_T_2907_addr] <= pages_T_2907_data;
    end
    if(pages_T_2911_en & pages_T_2911_mask) begin
      pages[pages_T_2911_addr] <= pages_T_2911_data;
    end
    if(pages_T_2915_en & pages_T_2915_mask) begin
      pages[pages_T_2915_addr] <= pages_T_2915_data;
    end
    if(reset) begin
      pageValid <= 6'h0;
    end else begin
      if(io_invalidate) begin
        pageValid <= {{5'd0}, 1'h0};
      end else begin
        if(r_btb_update_valid) begin
          if(doPageRepl) begin
            pageValid <= T_2916;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_581 == T_2550) begin
          useRAS_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_705 == T_2550) begin
          useRAS_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_784 == T_2550) begin
          useRAS_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_785 == T_2550) begin
          useRAS_3 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_786 == T_2550) begin
          useRAS_4 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_787 == T_2550) begin
          useRAS_5 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_788 == T_2550) begin
          useRAS_6 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_789 == T_2550) begin
          useRAS_7 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_790 == T_2550) begin
          useRAS_8 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_791 == T_2550) begin
          useRAS_9 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_792 == T_2550) begin
          useRAS_10 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_793 == T_2550) begin
          useRAS_11 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_794 == T_2550) begin
          useRAS_12 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_795 == T_2550) begin
          useRAS_13 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_796 == T_2550) begin
          useRAS_14 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_797 == T_2550) begin
          useRAS_15 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_798 == T_2550) begin
          useRAS_16 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_799 == T_2550) begin
          useRAS_17 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_800 == T_2550) begin
          useRAS_18 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_801 == T_2550) begin
          useRAS_19 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_802 == T_2550) begin
          useRAS_20 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_803 == T_2550) begin
          useRAS_21 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_804 == T_2550) begin
          useRAS_22 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_805 == T_2550) begin
          useRAS_23 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_806 == T_2550) begin
          useRAS_24 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_807 == T_2550) begin
          useRAS_25 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_808 == T_2550) begin
          useRAS_26 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_809 == T_2550) begin
          useRAS_27 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_810 == T_2550) begin
          useRAS_28 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_811 == T_2550) begin
          useRAS_29 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_812 == T_2550) begin
          useRAS_30 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_813 == T_2550) begin
          useRAS_31 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h20 == T_2550) begin
          useRAS_32 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h21 == T_2550) begin
          useRAS_33 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h22 == T_2550) begin
          useRAS_34 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h23 == T_2550) begin
          useRAS_35 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h24 == T_2550) begin
          useRAS_36 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h25 == T_2550) begin
          useRAS_37 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h26 == T_2550) begin
          useRAS_38 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h27 == T_2550) begin
          useRAS_39 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h28 == T_2550) begin
          useRAS_40 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h29 == T_2550) begin
          useRAS_41 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2a == T_2550) begin
          useRAS_42 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2b == T_2550) begin
          useRAS_43 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2c == T_2550) begin
          useRAS_44 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2d == T_2550) begin
          useRAS_45 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2e == T_2550) begin
          useRAS_46 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2f == T_2550) begin
          useRAS_47 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h30 == T_2550) begin
          useRAS_48 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h31 == T_2550) begin
          useRAS_49 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h32 == T_2550) begin
          useRAS_50 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h33 == T_2550) begin
          useRAS_51 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h34 == T_2550) begin
          useRAS_52 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h35 == T_2550) begin
          useRAS_53 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h36 == T_2550) begin
          useRAS_54 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h37 == T_2550) begin
          useRAS_55 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h38 == T_2550) begin
          useRAS_56 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h39 == T_2550) begin
          useRAS_57 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3a == T_2550) begin
          useRAS_58 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3b == T_2550) begin
          useRAS_59 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3c == T_2550) begin
          useRAS_60 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3d == T_2550) begin
          useRAS_61 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_581 == T_2550) begin
          isJump_0 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_705 == T_2550) begin
          isJump_1 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_784 == T_2550) begin
          isJump_2 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_785 == T_2550) begin
          isJump_3 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_786 == T_2550) begin
          isJump_4 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_787 == T_2550) begin
          isJump_5 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_788 == T_2550) begin
          isJump_6 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_789 == T_2550) begin
          isJump_7 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_790 == T_2550) begin
          isJump_8 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_791 == T_2550) begin
          isJump_9 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_792 == T_2550) begin
          isJump_10 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_793 == T_2550) begin
          isJump_11 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_794 == T_2550) begin
          isJump_12 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_795 == T_2550) begin
          isJump_13 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_796 == T_2550) begin
          isJump_14 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_797 == T_2550) begin
          isJump_15 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_798 == T_2550) begin
          isJump_16 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_799 == T_2550) begin
          isJump_17 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_800 == T_2550) begin
          isJump_18 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_801 == T_2550) begin
          isJump_19 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_802 == T_2550) begin
          isJump_20 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_803 == T_2550) begin
          isJump_21 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_804 == T_2550) begin
          isJump_22 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_805 == T_2550) begin
          isJump_23 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_806 == T_2550) begin
          isJump_24 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_807 == T_2550) begin
          isJump_25 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_808 == T_2550) begin
          isJump_26 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_809 == T_2550) begin
          isJump_27 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_810 == T_2550) begin
          isJump_28 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_811 == T_2550) begin
          isJump_29 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_812 == T_2550) begin
          isJump_30 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(GEN_813 == T_2550) begin
          isJump_31 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h20 == T_2550) begin
          isJump_32 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h21 == T_2550) begin
          isJump_33 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h22 == T_2550) begin
          isJump_34 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h23 == T_2550) begin
          isJump_35 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h24 == T_2550) begin
          isJump_36 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h25 == T_2550) begin
          isJump_37 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h26 == T_2550) begin
          isJump_38 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h27 == T_2550) begin
          isJump_39 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h28 == T_2550) begin
          isJump_40 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h29 == T_2550) begin
          isJump_41 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2a == T_2550) begin
          isJump_42 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2b == T_2550) begin
          isJump_43 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2c == T_2550) begin
          isJump_44 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2d == T_2550) begin
          isJump_45 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2e == T_2550) begin
          isJump_46 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2f == T_2550) begin
          isJump_47 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h30 == T_2550) begin
          isJump_48 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h31 == T_2550) begin
          isJump_49 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h32 == T_2550) begin
          isJump_50 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h33 == T_2550) begin
          isJump_51 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h34 == T_2550) begin
          isJump_52 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h35 == T_2550) begin
          isJump_53 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h36 == T_2550) begin
          isJump_54 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h37 == T_2550) begin
          isJump_55 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h38 == T_2550) begin
          isJump_56 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h39 == T_2550) begin
          isJump_57 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3a == T_2550) begin
          isJump_58 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3b == T_2550) begin
          isJump_59 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3c == T_2550) begin
          isJump_60 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3d == T_2550) begin
          isJump_61 <= GEN_1;
        end
      end
    end
    if(brIdx_T_2876_en & brIdx_T_2876_mask) begin
      brIdx[brIdx_T_2876_addr] <= brIdx_T_2876_data;
    end
    if(reset) begin
      T_1215 <= 1'h0;
    end else begin
      T_1215 <= io_btb_update_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_prediction_valid <= io_btb_update_bits_prediction_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_prediction_bits_taken <= io_btb_update_bits_prediction_bits_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_prediction_bits_mask <= io_btb_update_bits_prediction_bits_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_prediction_bits_bridx <= io_btb_update_bits_prediction_bits_bridx;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_prediction_bits_target <= io_btb_update_bits_prediction_bits_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_prediction_bits_entry <= io_btb_update_bits_prediction_bits_entry;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_prediction_bits_bht_history <= io_btb_update_bits_prediction_bits_bht_history;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_prediction_bits_bht_value <= io_btb_update_bits_prediction_bits_bht_value;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_pc <= io_btb_update_bits_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_target <= io_btb_update_bits_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_taken <= io_btb_update_bits_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_isJump <= io_btb_update_bits_isJump;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_isReturn <= io_btb_update_bits_isReturn;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_1216_br_pc <= io_btb_update_bits_br_pc;
      end
    end
    if(reset) begin
      nextRepl <= 6'h0;
    end else begin
      if(T_2482) begin
        if(T_2485) begin
          nextRepl <= {{5'd0}, 1'h0};
        end else begin
          nextRepl <= T_2488;
        end
      end
    end
    if(reset) begin
      T_2536 <= 3'h0;
    end else begin
      if(T_2534) begin
        if(T_2538) begin
          T_2536 <= {{2'd0}, 1'h0};
        end else begin
          T_2536 <= T_2541;
        end
      end
    end
    if(T_3616_T_3949_en & T_3616_T_3949_mask) begin
      T_3616[T_3616_T_3949_addr] <= T_3616_T_3949_data;
    end
    if(1'h0) begin
    end else begin
      if(T_3946) begin
        if(io_bht_update_bits_mispredict) begin
          T_3618 <= T_3960;
        end else begin
          if(T_3933) begin
            T_3618 <= T_3945;
          end
        end
      end else begin
        if(T_3933) begin
          T_3618 <= T_3945;
        end
      end
    end
    if(reset) begin
      T_3967 <= 2'h0;
    end else begin
      if(io_invalidate) begin
        T_3967 <= {{1'd0}, 1'h0};
      end else begin
        if(io_ras_update_valid) begin
          if(T_4311) begin
            if(T_4292) begin
              T_3967 <= T_4318;
            end else begin
              if(io_ras_update_bits_isCall) begin
                if(T_4295) begin
                  T_3967 <= T_4298;
                end
              end
            end
          end else begin
            if(io_ras_update_bits_isCall) begin
              if(T_4295) begin
                T_3967 <= T_4298;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_3969 <= 1'h0;
    end else begin
      if(io_ras_update_valid) begin
        if(T_4311) begin
          if(T_4292) begin
            T_3969 <= T_4325;
          end else begin
            if(io_ras_update_bits_isCall) begin
              T_3969 <= T_4305;
            end
          end
        end else begin
          if(io_ras_update_bits_isCall) begin
            T_3969 <= T_4305;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ras_update_valid) begin
        if(io_ras_update_bits_isCall) begin
          if(1'h0 == T_4305) begin
            T_3976_0 <= GEN_3;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ras_update_valid) begin
        if(io_ras_update_bits_isCall) begin
          if(T_4305) begin
            T_3976_1 <= GEN_3;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (r_btb_update_valid & T_2549) begin
          $fwrite(32'h80000002,"Assertion failed: BTB request != I$ target\n    at btb.scala:202 assert(io.req.bits.addr === r_btb_update.bits.target, \"BTB request != I$ target\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (r_btb_update_valid & T_2549) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (r_btb_update_valid & T_2549) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Queue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input  [63:0] io_enq_bits_datablock,
  input   io_deq_ready,
  output  io_deq_valid,
  output [31:0] io_deq_bits_data,
  output [63:0] io_deq_bits_datablock,
  output  io_count
);
  reg [31:0] ram_data [0:0];
  reg [31:0] GEN_0;
  wire [31:0] ram_data_T_744_data;
  wire  ram_data_T_744_addr;
  wire  ram_data_T_744_en;
  wire [31:0] ram_data_T_665_data;
  wire  ram_data_T_665_addr;
  wire  ram_data_T_665_mask;
  wire  ram_data_T_665_en;
  reg [63:0] ram_datablock [0:0];
  reg [63:0] GEN_1;
  wire [63:0] ram_datablock_T_744_data;
  wire  ram_datablock_T_744_addr;
  wire  ram_datablock_T_744_en;
  wire [63:0] ram_datablock_T_665_data;
  wire  ram_datablock_T_665_addr;
  wire  ram_datablock_T_665_mask;
  wire  ram_datablock_T_665_en;
  reg  maybe_full;
  reg [31:0] GEN_2;
  wire  T_662;
  wire  T_663;
  wire  do_enq;
  wire  T_664;
  wire  do_deq;
  wire  T_739;
  wire  GEN_7;
  wire  T_741;
  wire  GEN_8;
  wire [1:0] T_817;
  wire  ptr_diff;
  wire [1:0] T_819;
  assign io_enq_ready = GEN_8;
  assign io_deq_valid = T_741;
  assign io_deq_bits_data = ram_data_T_744_data;
  assign io_deq_bits_datablock = ram_datablock_T_744_data;
  assign io_count = T_819[0];
  assign ram_data_T_744_addr = 1'h0;
  assign ram_data_T_744_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_data_T_744_data = ram_data[ram_data_T_744_addr];
  `else
  assign ram_data_T_744_data = ram_data_T_744_addr >= 1'h1 ? $random : ram_data[ram_data_T_744_addr];
  `endif
  assign ram_data_T_665_data = io_enq_bits_data;
  assign ram_data_T_665_addr = 1'h0;
  assign ram_data_T_665_mask = do_enq;
  assign ram_data_T_665_en = do_enq;
  assign ram_datablock_T_744_addr = 1'h0;
  assign ram_datablock_T_744_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_datablock_T_744_data = ram_datablock[ram_datablock_T_744_addr];
  `else
  assign ram_datablock_T_744_data = ram_datablock_T_744_addr >= 1'h1 ? $random : ram_datablock[ram_datablock_T_744_addr];
  `endif
  assign ram_datablock_T_665_data = io_enq_bits_datablock;
  assign ram_datablock_T_665_addr = 1'h0;
  assign ram_datablock_T_665_mask = do_enq;
  assign ram_datablock_T_665_en = do_enq;
  assign T_662 = maybe_full == 1'h0;
  assign T_663 = io_enq_ready & io_enq_valid;
  assign do_enq = T_663;
  assign T_664 = io_deq_ready & io_deq_valid;
  assign do_deq = T_664;
  assign T_739 = do_enq != do_deq;
  assign GEN_7 = T_739 ? do_enq : maybe_full;
  assign T_741 = T_662 == 1'h0;
  assign GEN_8 = io_deq_ready ? 1'h1 : T_662;
  assign T_817 = 1'h0 - 1'h0;
  assign ptr_diff = T_817[0:0];
  assign T_819 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_0[31:0];
  GEN_1 = {2{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_datablock[initvar] = GEN_1[63:0];
  GEN_2 = {1{$random}};
  maybe_full = GEN_2[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_data_T_665_en & ram_data_T_665_mask) begin
      ram_data[ram_data_T_665_addr] <= ram_data_T_665_data;
    end
    if(ram_datablock_T_665_en & ram_datablock_T_665_mask) begin
      ram_datablock[ram_datablock_T_665_addr] <= ram_datablock_T_665_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_739) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Frontend(
  input   clk,
  input   reset,
  input   io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_pc,
  input   io_cpu_resp_ready,
  output  io_cpu_resp_valid,
  output [39:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data_0,
  output  io_cpu_resp_bits_mask,
  output  io_cpu_resp_bits_xcpt_if,
  output  io_cpu_btb_resp_valid,
  output  io_cpu_btb_resp_bits_taken,
  output  io_cpu_btb_resp_bits_mask,
  output  io_cpu_btb_resp_bits_bridx,
  output [38:0] io_cpu_btb_resp_bits_target,
  output [5:0] io_cpu_btb_resp_bits_entry,
  output [6:0] io_cpu_btb_resp_bits_bht_history,
  output [1:0] io_cpu_btb_resp_bits_bht_value,
  input   io_cpu_btb_update_valid,
  input   io_cpu_btb_update_bits_prediction_valid,
  input   io_cpu_btb_update_bits_prediction_bits_taken,
  input   io_cpu_btb_update_bits_prediction_bits_mask,
  input   io_cpu_btb_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_btb_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_btb_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
  input  [38:0] io_cpu_btb_update_bits_pc,
  input  [38:0] io_cpu_btb_update_bits_target,
  input   io_cpu_btb_update_bits_taken,
  input   io_cpu_btb_update_bits_isJump,
  input   io_cpu_btb_update_bits_isReturn,
  input  [38:0] io_cpu_btb_update_bits_br_pc,
  input   io_cpu_bht_update_valid,
  input   io_cpu_bht_update_bits_prediction_valid,
  input   io_cpu_bht_update_bits_prediction_bits_taken,
  input   io_cpu_bht_update_bits_prediction_bits_mask,
  input   io_cpu_bht_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_bht_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_bht_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_bht_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
  input  [38:0] io_cpu_bht_update_bits_pc,
  input   io_cpu_bht_update_bits_taken,
  input   io_cpu_bht_update_bits_mispredict,
  input   io_cpu_ras_update_valid,
  input   io_cpu_ras_update_bits_isCall,
  input   io_cpu_ras_update_bits_isReturn,
  input  [38:0] io_cpu_ras_update_bits_returnAddr,
  input   io_cpu_ras_update_bits_prediction_valid,
  input   io_cpu_ras_update_bits_prediction_bits_taken,
  input   io_cpu_ras_update_bits_prediction_bits_mask,
  input   io_cpu_ras_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_ras_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_ras_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_ras_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
  input   io_cpu_flush_icache,
  input   io_cpu_flush_tlb,
  output [39:0] io_cpu_npc,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_addr,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [19:0] io_ptw_resp_bits_pte_ppn,
  input  [2:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_r,
  input  [3:0] io_ptw_resp_bits_pte_typ,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [4:0] io_ptw_status_zero1,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_req_valid;
  wire [38:0] icache_io_req_bits_addr;
  wire [19:0] icache_io_s1_ppn;
  wire  icache_io_s1_kill;
  wire  icache_io_resp_ready;
  wire  icache_io_resp_valid;
  wire [31:0] icache_io_resp_bits_data;
  wire [63:0] icache_io_resp_bits_datablock;
  wire  icache_io_invalidate;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire [1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [11:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire [1:0] icache_io_mem_grant_bits_client_xact_id;
  wire [2:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  tlb_clk;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [27:0] tlb_io_req_bits_vpn;
  wire  tlb_io_req_bits_passthrough;
  wire  tlb_io_req_bits_instruction;
  wire  tlb_io_req_bits_store;
  wire  tlb_io_resp_miss;
  wire [19:0] tlb_io_resp_ppn;
  wire  tlb_io_resp_xcpt_ld;
  wire  tlb_io_resp_xcpt_st;
  wire  tlb_io_resp_xcpt_if;
  wire [7:0] tlb_io_resp_hit_idx;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [26:0] tlb_io_ptw_req_bits_addr;
  wire [1:0] tlb_io_ptw_req_bits_prv;
  wire  tlb_io_ptw_req_bits_store;
  wire  tlb_io_ptw_req_bits_fetch;
  wire  tlb_io_ptw_resp_valid;
  wire [19:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire [2:0] tlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire [3:0] tlb_io_ptw_resp_bits_pte_typ;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire [6:0] tlb_io_ptw_ptbr_asid;
  wire [37:0] tlb_io_ptw_ptbr_ppn;
  wire  tlb_io_ptw_invalidate;
  wire  tlb_io_ptw_status_debug;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_sd;
  wire [30:0] tlb_io_ptw_status_zero3;
  wire  tlb_io_ptw_status_sd_rv32;
  wire [1:0] tlb_io_ptw_status_zero2;
  wire [4:0] tlb_io_ptw_status_vm;
  wire [4:0] tlb_io_ptw_status_zero1;
  wire  tlb_io_ptw_status_pum;
  wire  tlb_io_ptw_status_mprv;
  wire [1:0] tlb_io_ptw_status_xs;
  wire [1:0] tlb_io_ptw_status_fs;
  wire [1:0] tlb_io_ptw_status_mpp;
  wire [1:0] tlb_io_ptw_status_hpp;
  wire  tlb_io_ptw_status_spp;
  wire  tlb_io_ptw_status_mpie;
  wire  tlb_io_ptw_status_hpie;
  wire  tlb_io_ptw_status_spie;
  wire  tlb_io_ptw_status_upie;
  wire  tlb_io_ptw_status_mie;
  wire  tlb_io_ptw_status_hie;
  wire  tlb_io_ptw_status_sie;
  wire  tlb_io_ptw_status_uie;
  reg [39:0] s1_pc_;
  reg [63:0] GEN_10;
  wire [39:0] T_1302;
  wire [39:0] GEN_21;
  wire [39:0] T_1304;
  wire [39:0] s1_pc;
  reg  s1_same_block;
  reg [31:0] GEN_22;
  reg  s2_valid;
  reg [31:0] GEN_28;
  reg [39:0] s2_pc;
  reg [63:0] GEN_29;
  reg  s2_btb_resp_valid;
  reg [31:0] GEN_30;
  reg  s2_btb_resp_bits_taken;
  reg [31:0] GEN_31;
  reg  s2_btb_resp_bits_mask;
  reg [31:0] GEN_32;
  reg  s2_btb_resp_bits_bridx;
  reg [31:0] GEN_33;
  reg [38:0] s2_btb_resp_bits_target;
  reg [63:0] GEN_34;
  reg [5:0] s2_btb_resp_bits_entry;
  reg [31:0] GEN_35;
  reg [6:0] s2_btb_resp_bits_bht_history;
  reg [31:0] GEN_36;
  reg [1:0] s2_btb_resp_bits_bht_value;
  reg [31:0] GEN_37;
  reg  s2_xcpt_if;
  reg [31:0] GEN_38;
  wire  s2_resp_valid;
  wire [63:0] s2_resp_data;
  wire [39:0] T_1329;
  wire [39:0] T_1331;
  wire [39:0] T_1332;
  wire [39:0] GEN_23;
  wire [40:0] T_1334;
  wire [39:0] ntpc_0;
  wire  T_1335;
  wire  T_1336;
  wire  T_1337;
  wire [40:0] ntpc;
  wire [40:0] predicted_npc;
  wire  T_1339;
  wire  icmiss;
  wire [40:0] npc;
  wire  T_1341;
  wire  T_1343;
  wire  T_1344;
  wire [40:0] GEN_24;
  wire [40:0] T_1346;
  wire [39:0] GEN_25;
  wire [39:0] T_1348;
  wire [40:0] GEN_26;
  wire  T_1349;
  wire  T_1350;
  wire  s0_same_block;
  wire  T_1352;
  wire  stall;
  wire  T_1354;
  wire  T_1356;
  wire  T_1357;
  wire [39:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire [40:0] GEN_3;
  wire  GEN_4;
  wire [39:0] GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [40:0] GEN_8;
  wire  GEN_9;
  wire  BTB_1_clk;
  wire  BTB_1_reset;
  wire  BTB_1_io_req_valid;
  wire [38:0] BTB_1_io_req_bits_addr;
  wire  BTB_1_io_resp_valid;
  wire  BTB_1_io_resp_bits_taken;
  wire  BTB_1_io_resp_bits_mask;
  wire  BTB_1_io_resp_bits_bridx;
  wire [38:0] BTB_1_io_resp_bits_target;
  wire [5:0] BTB_1_io_resp_bits_entry;
  wire [6:0] BTB_1_io_resp_bits_bht_history;
  wire [1:0] BTB_1_io_resp_bits_bht_value;
  wire  BTB_1_io_btb_update_valid;
  wire  BTB_1_io_btb_update_bits_prediction_valid;
  wire  BTB_1_io_btb_update_bits_prediction_bits_taken;
  wire  BTB_1_io_btb_update_bits_prediction_bits_mask;
  wire  BTB_1_io_btb_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1_io_btb_update_bits_prediction_bits_target;
  wire [5:0] BTB_1_io_btb_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1_io_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1_io_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] BTB_1_io_btb_update_bits_pc;
  wire [38:0] BTB_1_io_btb_update_bits_target;
  wire  BTB_1_io_btb_update_bits_taken;
  wire  BTB_1_io_btb_update_bits_isJump;
  wire  BTB_1_io_btb_update_bits_isReturn;
  wire [38:0] BTB_1_io_btb_update_bits_br_pc;
  wire  BTB_1_io_bht_update_valid;
  wire  BTB_1_io_bht_update_bits_prediction_valid;
  wire  BTB_1_io_bht_update_bits_prediction_bits_taken;
  wire  BTB_1_io_bht_update_bits_prediction_bits_mask;
  wire  BTB_1_io_bht_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1_io_bht_update_bits_prediction_bits_target;
  wire [5:0] BTB_1_io_bht_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1_io_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1_io_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] BTB_1_io_bht_update_bits_pc;
  wire  BTB_1_io_bht_update_bits_taken;
  wire  BTB_1_io_bht_update_bits_mispredict;
  wire  BTB_1_io_ras_update_valid;
  wire  BTB_1_io_ras_update_bits_isCall;
  wire  BTB_1_io_ras_update_bits_isReturn;
  wire [38:0] BTB_1_io_ras_update_bits_returnAddr;
  wire  BTB_1_io_ras_update_bits_prediction_valid;
  wire  BTB_1_io_ras_update_bits_prediction_bits_taken;
  wire  BTB_1_io_ras_update_bits_prediction_bits_mask;
  wire  BTB_1_io_ras_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1_io_ras_update_bits_prediction_bits_target;
  wire [5:0] BTB_1_io_ras_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1_io_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1_io_ras_update_bits_prediction_bits_bht_value;
  wire  BTB_1_io_invalidate;
  wire  T_1370;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [38:0] GEN_15;
  wire [5:0] GEN_16;
  wire [6:0] GEN_17;
  wire [1:0] GEN_18;
  wire  T_1372;
  wire [39:0] T_1373;
  wire [40:0] GEN_19;
  wire  GEN_20;
  wire [27:0] T_1380;
  wire  T_1387;
  wire  T_1388;
  wire  T_1389;
  wire  T_1390;
  wire  T_1391;
  wire  T_1392;
  wire  T_1393;
  wire  T_1394;
  wire [40:0] T_1395;
  wire  Queue_1_clk;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [31:0] Queue_1_io_enq_bits_data;
  wire [63:0] Queue_1_io_enq_bits_datablock;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [31:0] Queue_1_io_deq_bits_data;
  wire [63:0] Queue_1_io_deq_bits_datablock;
  wire  Queue_1_io_count;
  wire  T_1471;
  wire  T_1472;
  wire  T_1473;
  wire [5:0] GEN_27;
  wire [5:0] T_1474;
  wire [63:0] fetch_data;
  wire [31:0] T_1475;
  ICache icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_ppn(icache_io_s1_ppn),
    .io_s1_kill(icache_io_s1_kill),
    .io_resp_ready(icache_io_resp_ready),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_datablock(icache_io_resp_bits_datablock),
    .io_invalidate(icache_io_invalidate),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  TLB tlb (
    .clk(tlb_clk),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vpn(tlb_io_req_bits_vpn),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_store(tlb_io_req_bits_store),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_ppn(tlb_io_resp_ppn),
    .io_resp_xcpt_ld(tlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(tlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(tlb_io_resp_xcpt_if),
    .io_resp_hit_idx(tlb_io_resp_hit_idx),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_prv(tlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_store(tlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(tlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(tlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_typ(tlb_io_ptw_resp_bits_pte_typ),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(tlb_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(tlb_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(tlb_io_ptw_invalidate),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_sd(tlb_io_ptw_status_sd),
    .io_ptw_status_zero3(tlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(tlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(tlb_io_ptw_status_zero2),
    .io_ptw_status_vm(tlb_io_ptw_status_vm),
    .io_ptw_status_zero1(tlb_io_ptw_status_zero1),
    .io_ptw_status_pum(tlb_io_ptw_status_pum),
    .io_ptw_status_mprv(tlb_io_ptw_status_mprv),
    .io_ptw_status_xs(tlb_io_ptw_status_xs),
    .io_ptw_status_fs(tlb_io_ptw_status_fs),
    .io_ptw_status_mpp(tlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(tlb_io_ptw_status_hpp),
    .io_ptw_status_spp(tlb_io_ptw_status_spp),
    .io_ptw_status_mpie(tlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(tlb_io_ptw_status_hpie),
    .io_ptw_status_spie(tlb_io_ptw_status_spie),
    .io_ptw_status_upie(tlb_io_ptw_status_upie),
    .io_ptw_status_mie(tlb_io_ptw_status_mie),
    .io_ptw_status_hie(tlb_io_ptw_status_hie),
    .io_ptw_status_sie(tlb_io_ptw_status_sie),
    .io_ptw_status_uie(tlb_io_ptw_status_uie)
  );
  BTB BTB_1 (
    .clk(BTB_1_clk),
    .reset(BTB_1_reset),
    .io_req_valid(BTB_1_io_req_valid),
    .io_req_bits_addr(BTB_1_io_req_bits_addr),
    .io_resp_valid(BTB_1_io_resp_valid),
    .io_resp_bits_taken(BTB_1_io_resp_bits_taken),
    .io_resp_bits_mask(BTB_1_io_resp_bits_mask),
    .io_resp_bits_bridx(BTB_1_io_resp_bits_bridx),
    .io_resp_bits_target(BTB_1_io_resp_bits_target),
    .io_resp_bits_entry(BTB_1_io_resp_bits_entry),
    .io_resp_bits_bht_history(BTB_1_io_resp_bits_bht_history),
    .io_resp_bits_bht_value(BTB_1_io_resp_bits_bht_value),
    .io_btb_update_valid(BTB_1_io_btb_update_valid),
    .io_btb_update_bits_prediction_valid(BTB_1_io_btb_update_bits_prediction_valid),
    .io_btb_update_bits_prediction_bits_taken(BTB_1_io_btb_update_bits_prediction_bits_taken),
    .io_btb_update_bits_prediction_bits_mask(BTB_1_io_btb_update_bits_prediction_bits_mask),
    .io_btb_update_bits_prediction_bits_bridx(BTB_1_io_btb_update_bits_prediction_bits_bridx),
    .io_btb_update_bits_prediction_bits_target(BTB_1_io_btb_update_bits_prediction_bits_target),
    .io_btb_update_bits_prediction_bits_entry(BTB_1_io_btb_update_bits_prediction_bits_entry),
    .io_btb_update_bits_prediction_bits_bht_history(BTB_1_io_btb_update_bits_prediction_bits_bht_history),
    .io_btb_update_bits_prediction_bits_bht_value(BTB_1_io_btb_update_bits_prediction_bits_bht_value),
    .io_btb_update_bits_pc(BTB_1_io_btb_update_bits_pc),
    .io_btb_update_bits_target(BTB_1_io_btb_update_bits_target),
    .io_btb_update_bits_taken(BTB_1_io_btb_update_bits_taken),
    .io_btb_update_bits_isJump(BTB_1_io_btb_update_bits_isJump),
    .io_btb_update_bits_isReturn(BTB_1_io_btb_update_bits_isReturn),
    .io_btb_update_bits_br_pc(BTB_1_io_btb_update_bits_br_pc),
    .io_bht_update_valid(BTB_1_io_bht_update_valid),
    .io_bht_update_bits_prediction_valid(BTB_1_io_bht_update_bits_prediction_valid),
    .io_bht_update_bits_prediction_bits_taken(BTB_1_io_bht_update_bits_prediction_bits_taken),
    .io_bht_update_bits_prediction_bits_mask(BTB_1_io_bht_update_bits_prediction_bits_mask),
    .io_bht_update_bits_prediction_bits_bridx(BTB_1_io_bht_update_bits_prediction_bits_bridx),
    .io_bht_update_bits_prediction_bits_target(BTB_1_io_bht_update_bits_prediction_bits_target),
    .io_bht_update_bits_prediction_bits_entry(BTB_1_io_bht_update_bits_prediction_bits_entry),
    .io_bht_update_bits_prediction_bits_bht_history(BTB_1_io_bht_update_bits_prediction_bits_bht_history),
    .io_bht_update_bits_prediction_bits_bht_value(BTB_1_io_bht_update_bits_prediction_bits_bht_value),
    .io_bht_update_bits_pc(BTB_1_io_bht_update_bits_pc),
    .io_bht_update_bits_taken(BTB_1_io_bht_update_bits_taken),
    .io_bht_update_bits_mispredict(BTB_1_io_bht_update_bits_mispredict),
    .io_ras_update_valid(BTB_1_io_ras_update_valid),
    .io_ras_update_bits_isCall(BTB_1_io_ras_update_bits_isCall),
    .io_ras_update_bits_isReturn(BTB_1_io_ras_update_bits_isReturn),
    .io_ras_update_bits_returnAddr(BTB_1_io_ras_update_bits_returnAddr),
    .io_ras_update_bits_prediction_valid(BTB_1_io_ras_update_bits_prediction_valid),
    .io_ras_update_bits_prediction_bits_taken(BTB_1_io_ras_update_bits_prediction_bits_taken),
    .io_ras_update_bits_prediction_bits_mask(BTB_1_io_ras_update_bits_prediction_bits_mask),
    .io_ras_update_bits_prediction_bits_bridx(BTB_1_io_ras_update_bits_prediction_bits_bridx),
    .io_ras_update_bits_prediction_bits_target(BTB_1_io_ras_update_bits_prediction_bits_target),
    .io_ras_update_bits_prediction_bits_entry(BTB_1_io_ras_update_bits_prediction_bits_entry),
    .io_ras_update_bits_prediction_bits_bht_history(BTB_1_io_ras_update_bits_prediction_bits_bht_history),
    .io_ras_update_bits_prediction_bits_bht_value(BTB_1_io_ras_update_bits_prediction_bits_bht_value),
    .io_invalidate(BTB_1_io_invalidate)
  );
  Queue Queue_1 (
    .clk(Queue_1_clk),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_datablock(Queue_1_io_enq_bits_datablock),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_datablock(Queue_1_io_deq_bits_datablock),
    .io_count(Queue_1_io_count)
  );
  assign io_cpu_resp_valid = T_1394;
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_bits_data_0 = T_1475;
  assign io_cpu_resp_bits_mask = 1'h1;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_bits_mask = s2_btb_resp_bits_mask;
  assign io_cpu_btb_resp_bits_bridx = s2_btb_resp_bits_bridx;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign io_cpu_npc = T_1395[39:0];
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_req_valid = T_1388;
  assign icache_io_req_bits_addr = io_cpu_npc[38:0];
  assign icache_io_s1_ppn = tlb_io_resp_ppn;
  assign icache_io_s1_kill = T_1392;
  assign icache_io_resp_ready = Queue_1_io_enq_ready;
  assign icache_io_invalidate = io_cpu_flush_icache;
  assign icache_io_mem_acquire_ready = io_mem_acquire_ready;
  assign icache_io_mem_grant_valid = io_mem_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign tlb_clk = clk;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = T_1370;
  assign tlb_io_req_bits_vpn = T_1380;
  assign tlb_io_req_bits_passthrough = 1'h0;
  assign tlb_io_req_bits_instruction = 1'h1;
  assign tlb_io_req_bits_store = 1'h0;
  assign tlb_io_ptw_req_ready = io_ptw_req_ready;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign tlb_io_ptw_resp_bits_pte_typ = io_ptw_resp_bits_pte_typ;
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign tlb_io_ptw_ptbr_asid = io_ptw_ptbr_asid;
  assign tlb_io_ptw_ptbr_ppn = io_ptw_ptbr_ppn;
  assign tlb_io_ptw_invalidate = io_ptw_invalidate;
  assign tlb_io_ptw_status_debug = io_ptw_status_debug;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_sd = io_ptw_status_sd;
  assign tlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign tlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign tlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign tlb_io_ptw_status_vm = io_ptw_status_vm;
  assign tlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign tlb_io_ptw_status_pum = io_ptw_status_pum;
  assign tlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign tlb_io_ptw_status_xs = io_ptw_status_xs;
  assign tlb_io_ptw_status_fs = io_ptw_status_fs;
  assign tlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign tlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign tlb_io_ptw_status_spp = io_ptw_status_spp;
  assign tlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign tlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign tlb_io_ptw_status_spie = io_ptw_status_spie;
  assign tlb_io_ptw_status_upie = io_ptw_status_upie;
  assign tlb_io_ptw_status_mie = io_ptw_status_mie;
  assign tlb_io_ptw_status_hie = io_ptw_status_hie;
  assign tlb_io_ptw_status_sie = io_ptw_status_sie;
  assign tlb_io_ptw_status_uie = io_ptw_status_uie;
  assign T_1302 = ~ s1_pc_;
  assign GEN_21 = {{38'd0}, 2'h3};
  assign T_1304 = T_1302 | GEN_21;
  assign s1_pc = ~ T_1304;
  assign s2_resp_valid = Queue_1_io_deq_valid;
  assign s2_resp_data = Queue_1_io_deq_bits_datablock;
  assign T_1329 = ~ s1_pc;
  assign T_1331 = T_1329 | GEN_21;
  assign T_1332 = ~ T_1331;
  assign GEN_23 = {{37'd0}, 3'h4};
  assign T_1334 = T_1332 + GEN_23;
  assign ntpc_0 = T_1334[39:0];
  assign T_1335 = s1_pc[38];
  assign T_1336 = ntpc_0[38];
  assign T_1337 = T_1335 & T_1336;
  assign ntpc = {T_1337,ntpc_0};
  assign predicted_npc = GEN_19;
  assign T_1339 = s2_resp_valid == 1'h0;
  assign icmiss = s2_valid & T_1339;
  assign npc = icmiss ? {{1'd0}, s2_pc} : predicted_npc;
  assign T_1341 = icmiss == 1'h0;
  assign T_1343 = io_cpu_req_valid == 1'h0;
  assign T_1344 = T_1341 & T_1343;
  assign GEN_24 = {{37'd0}, 4'h8};
  assign T_1346 = ntpc & GEN_24;
  assign GEN_25 = {{36'd0}, 4'h8};
  assign T_1348 = s1_pc & GEN_25;
  assign GEN_26 = {{1'd0}, T_1348};
  assign T_1349 = T_1346 == GEN_26;
  assign T_1350 = T_1344 & T_1349;
  assign s0_same_block = GEN_20;
  assign T_1352 = io_cpu_resp_ready == 1'h0;
  assign stall = io_cpu_resp_valid & T_1352;
  assign T_1354 = stall == 1'h0;
  assign T_1356 = tlb_io_resp_miss == 1'h0;
  assign T_1357 = s0_same_block & T_1356;
  assign GEN_0 = T_1341 ? s1_pc : s2_pc;
  assign GEN_1 = T_1341 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign GEN_2 = T_1354 ? T_1357 : s1_same_block;
  assign GEN_3 = T_1354 ? npc : {{1'd0}, s1_pc_};
  assign GEN_4 = T_1354 ? T_1341 : s2_valid;
  assign GEN_5 = T_1354 ? GEN_0 : s2_pc;
  assign GEN_6 = T_1354 ? GEN_1 : s2_xcpt_if;
  assign GEN_7 = io_cpu_req_valid ? 1'h0 : GEN_2;
  assign GEN_8 = io_cpu_req_valid ? {{1'd0}, io_cpu_req_bits_pc} : GEN_3;
  assign GEN_9 = io_cpu_req_valid ? 1'h0 : GEN_4;
  assign BTB_1_clk = clk;
  assign BTB_1_reset = reset;
  assign BTB_1_io_req_valid = T_1370;
  assign BTB_1_io_req_bits_addr = s1_pc[38:0];
  assign BTB_1_io_btb_update_valid = io_cpu_btb_update_valid;
  assign BTB_1_io_btb_update_bits_prediction_valid = io_cpu_btb_update_bits_prediction_valid;
  assign BTB_1_io_btb_update_bits_prediction_bits_taken = io_cpu_btb_update_bits_prediction_bits_taken;
  assign BTB_1_io_btb_update_bits_prediction_bits_mask = io_cpu_btb_update_bits_prediction_bits_mask;
  assign BTB_1_io_btb_update_bits_prediction_bits_bridx = io_cpu_btb_update_bits_prediction_bits_bridx;
  assign BTB_1_io_btb_update_bits_prediction_bits_target = io_cpu_btb_update_bits_prediction_bits_target;
  assign BTB_1_io_btb_update_bits_prediction_bits_entry = io_cpu_btb_update_bits_prediction_bits_entry;
  assign BTB_1_io_btb_update_bits_prediction_bits_bht_history = io_cpu_btb_update_bits_prediction_bits_bht_history;
  assign BTB_1_io_btb_update_bits_prediction_bits_bht_value = io_cpu_btb_update_bits_prediction_bits_bht_value;
  assign BTB_1_io_btb_update_bits_pc = io_cpu_btb_update_bits_pc;
  assign BTB_1_io_btb_update_bits_target = io_cpu_btb_update_bits_target;
  assign BTB_1_io_btb_update_bits_taken = io_cpu_btb_update_bits_taken;
  assign BTB_1_io_btb_update_bits_isJump = io_cpu_btb_update_bits_isJump;
  assign BTB_1_io_btb_update_bits_isReturn = io_cpu_btb_update_bits_isReturn;
  assign BTB_1_io_btb_update_bits_br_pc = io_cpu_btb_update_bits_br_pc;
  assign BTB_1_io_bht_update_valid = io_cpu_bht_update_valid;
  assign BTB_1_io_bht_update_bits_prediction_valid = io_cpu_bht_update_bits_prediction_valid;
  assign BTB_1_io_bht_update_bits_prediction_bits_taken = io_cpu_bht_update_bits_prediction_bits_taken;
  assign BTB_1_io_bht_update_bits_prediction_bits_mask = io_cpu_bht_update_bits_prediction_bits_mask;
  assign BTB_1_io_bht_update_bits_prediction_bits_bridx = io_cpu_bht_update_bits_prediction_bits_bridx;
  assign BTB_1_io_bht_update_bits_prediction_bits_target = io_cpu_bht_update_bits_prediction_bits_target;
  assign BTB_1_io_bht_update_bits_prediction_bits_entry = io_cpu_bht_update_bits_prediction_bits_entry;
  assign BTB_1_io_bht_update_bits_prediction_bits_bht_history = io_cpu_bht_update_bits_prediction_bits_bht_history;
  assign BTB_1_io_bht_update_bits_prediction_bits_bht_value = io_cpu_bht_update_bits_prediction_bits_bht_value;
  assign BTB_1_io_bht_update_bits_pc = io_cpu_bht_update_bits_pc;
  assign BTB_1_io_bht_update_bits_taken = io_cpu_bht_update_bits_taken;
  assign BTB_1_io_bht_update_bits_mispredict = io_cpu_bht_update_bits_mispredict;
  assign BTB_1_io_ras_update_valid = io_cpu_ras_update_valid;
  assign BTB_1_io_ras_update_bits_isCall = io_cpu_ras_update_bits_isCall;
  assign BTB_1_io_ras_update_bits_isReturn = io_cpu_ras_update_bits_isReturn;
  assign BTB_1_io_ras_update_bits_returnAddr = io_cpu_ras_update_bits_returnAddr;
  assign BTB_1_io_ras_update_bits_prediction_valid = io_cpu_ras_update_bits_prediction_valid;
  assign BTB_1_io_ras_update_bits_prediction_bits_taken = io_cpu_ras_update_bits_prediction_bits_taken;
  assign BTB_1_io_ras_update_bits_prediction_bits_mask = io_cpu_ras_update_bits_prediction_bits_mask;
  assign BTB_1_io_ras_update_bits_prediction_bits_bridx = io_cpu_ras_update_bits_prediction_bits_bridx;
  assign BTB_1_io_ras_update_bits_prediction_bits_target = io_cpu_ras_update_bits_prediction_bits_target;
  assign BTB_1_io_ras_update_bits_prediction_bits_entry = io_cpu_ras_update_bits_prediction_bits_entry;
  assign BTB_1_io_ras_update_bits_prediction_bits_bht_history = io_cpu_ras_update_bits_prediction_bits_bht_history;
  assign BTB_1_io_ras_update_bits_prediction_bits_bht_value = io_cpu_ras_update_bits_prediction_bits_bht_value;
  assign BTB_1_io_invalidate = 1'h0;
  assign T_1370 = T_1354 & T_1341;
  assign GEN_11 = T_1370 ? BTB_1_io_resp_valid : s2_btb_resp_valid;
  assign GEN_12 = T_1370 ? BTB_1_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign GEN_13 = T_1370 ? BTB_1_io_resp_bits_mask : s2_btb_resp_bits_mask;
  assign GEN_14 = T_1370 ? BTB_1_io_resp_bits_bridx : s2_btb_resp_bits_bridx;
  assign GEN_15 = T_1370 ? BTB_1_io_resp_bits_target : s2_btb_resp_bits_target;
  assign GEN_16 = T_1370 ? BTB_1_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign GEN_17 = T_1370 ? BTB_1_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign GEN_18 = T_1370 ? BTB_1_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T_1372 = BTB_1_io_resp_bits_target[38];
  assign T_1373 = {T_1372,BTB_1_io_resp_bits_target};
  assign GEN_19 = BTB_1_io_resp_bits_taken ? {{1'd0}, T_1373} : ntpc;
  assign GEN_20 = BTB_1_io_resp_bits_taken ? 1'h0 : T_1350;
  assign T_1380 = s1_pc[39:12];
  assign T_1387 = s0_same_block == 1'h0;
  assign T_1388 = T_1354 & T_1387;
  assign T_1389 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T_1390 = T_1389 | tlb_io_resp_xcpt_if;
  assign T_1391 = T_1390 | icmiss;
  assign T_1392 = T_1391 | io_cpu_flush_tlb;
  assign T_1393 = s2_xcpt_if | s2_resp_valid;
  assign T_1394 = s2_valid & T_1393;
  assign T_1395 = io_cpu_req_valid ? {{1'd0}, io_cpu_req_bits_pc} : npc;
  assign Queue_1_clk = clk;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = icache_io_resp_valid;
  assign Queue_1_io_enq_bits_data = icache_io_resp_bits_data;
  assign Queue_1_io_enq_bits_datablock = icache_io_resp_bits_datablock;
  assign Queue_1_io_deq_ready = T_1472;
  assign T_1471 = s1_same_block == 1'h0;
  assign T_1472 = T_1354 & T_1471;
  assign T_1473 = s2_pc[2];
  assign GEN_27 = {{5'd0}, T_1473};
  assign T_1474 = GEN_27 << 5;
  assign fetch_data = s2_resp_data >> T_1474;
  assign T_1475 = fetch_data[31:0];
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_10 = {2{$random}};
  s1_pc_ = GEN_10[39:0];
  GEN_22 = {1{$random}};
  s1_same_block = GEN_22[0:0];
  GEN_28 = {1{$random}};
  s2_valid = GEN_28[0:0];
  GEN_29 = {2{$random}};
  s2_pc = GEN_29[39:0];
  GEN_30 = {1{$random}};
  s2_btb_resp_valid = GEN_30[0:0];
  GEN_31 = {1{$random}};
  s2_btb_resp_bits_taken = GEN_31[0:0];
  GEN_32 = {1{$random}};
  s2_btb_resp_bits_mask = GEN_32[0:0];
  GEN_33 = {1{$random}};
  s2_btb_resp_bits_bridx = GEN_33[0:0];
  GEN_34 = {2{$random}};
  s2_btb_resp_bits_target = GEN_34[38:0];
  GEN_35 = {1{$random}};
  s2_btb_resp_bits_entry = GEN_35[5:0];
  GEN_36 = {1{$random}};
  s2_btb_resp_bits_bht_history = GEN_36[6:0];
  GEN_37 = {1{$random}};
  s2_btb_resp_bits_bht_value = GEN_37[1:0];
  GEN_38 = {1{$random}};
  s2_xcpt_if = GEN_38[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      s1_pc_ <= GEN_8[39:0];
    end
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_same_block <= 1'h0;
      end else begin
        if(T_1354) begin
          s1_same_block <= T_1357;
        end
      end
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else begin
      if(io_cpu_req_valid) begin
        s2_valid <= 1'h0;
      end else begin
        if(T_1354) begin
          s2_valid <= T_1341;
        end
      end
    end
    if(reset) begin
      s2_pc <= {{27'd0}, 13'h1000};
    end else begin
      if(T_1354) begin
        if(T_1341) begin
          s2_pc <= s1_pc;
        end
      end
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else begin
      if(T_1370) begin
        s2_btb_resp_valid <= BTB_1_io_resp_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1370) begin
        s2_btb_resp_bits_taken <= BTB_1_io_resp_bits_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1370) begin
        s2_btb_resp_bits_mask <= BTB_1_io_resp_bits_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1370) begin
        s2_btb_resp_bits_bridx <= BTB_1_io_resp_bits_bridx;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1370) begin
        s2_btb_resp_bits_target <= BTB_1_io_resp_bits_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1370) begin
        s2_btb_resp_bits_entry <= BTB_1_io_resp_bits_entry;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1370) begin
        s2_btb_resp_bits_bht_history <= BTB_1_io_resp_bits_bht_history;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1370) begin
        s2_btb_resp_bits_bht_value <= BTB_1_io_resp_bits_bht_value;
      end
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else begin
      if(T_1354) begin
        if(T_1341) begin
          s2_xcpt_if <= tlb_io_resp_xcpt_if;
        end
      end
    end
  end
endmodule
module WritebackUnit(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [2:0] io_req_bits_addr_beat,
  input  [25:0] io_req_bits_addr_block,
  input  [1:0] io_req_bits_client_xact_id,
  input   io_req_bits_voluntary,
  input  [2:0] io_req_bits_r_type,
  input  [63:0] io_req_bits_data,
  input  [3:0] io_req_bits_way_en,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_data_req_ready,
  output  io_data_req_valid,
  output [3:0] io_data_req_bits_way_en,
  output [11:0] io_data_req_bits_addr,
  input  [63:0] io_data_resp,
  input   io_release_ready,
  output  io_release_valid,
  output [2:0] io_release_bits_addr_beat,
  output [25:0] io_release_bits_addr_block,
  output [1:0] io_release_bits_client_xact_id,
  output  io_release_bits_voluntary,
  output [2:0] io_release_bits_r_type,
  output [63:0] io_release_bits_data
);
  reg  active;
  reg [31:0] GEN_6;
  reg  r1_data_req_fired;
  reg [31:0] GEN_7;
  reg  r2_data_req_fired;
  reg [31:0] GEN_8;
  reg [3:0] data_req_cnt;
  reg [31:0] GEN_10;
  wire  T_748;
  reg [2:0] beat_cnt;
  reg [31:0] GEN_33;
  wire [2:0] GEN_29;
  wire [3:0] T_753;
  wire [2:0] T_754;
  wire [2:0] GEN_0;
  reg [2:0] req_addr_beat;
  reg [31:0] GEN_34;
  reg [25:0] req_addr_block;
  reg [31:0] GEN_35;
  reg [1:0] req_client_xact_id;
  reg [31:0] GEN_36;
  reg  req_voluntary;
  reg [31:0] GEN_37;
  reg [2:0] req_r_type;
  reg [31:0] GEN_38;
  reg [63:0] req_data;
  reg [63:0] GEN_39;
  reg [3:0] req_way_en;
  reg [31:0] GEN_40;
  wire  T_864;
  wire  T_865;
  wire  T_866;
  wire [3:0] GEN_30;
  wire [4:0] T_869;
  wire [3:0] T_870;
  wire [3:0] GEN_2;
  wire  T_872;
  wire [1:0] T_879;
  wire [3:0] GEN_31;
  wire [4:0] T_880;
  wire [3:0] T_881;
  wire  GEN_3;
  wire  GEN_4;
  wire [3:0] GEN_5;
  wire  T_885;
  wire  T_887;
  wire  T_890;
  wire  GEN_9;
  wire  GEN_11;
  wire  GEN_12;
  wire [3:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [3:0] GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  T_891;
  wire  GEN_20;
  wire [3:0] GEN_21;
  wire [2:0] GEN_22;
  wire [25:0] GEN_23;
  wire [1:0] GEN_24;
  wire  GEN_25;
  wire [2:0] GEN_26;
  wire [63:0] GEN_27;
  wire [3:0] GEN_28;
  wire  T_895;
  wire [5:0] req_idx;
  wire  fire;
  wire [19:0] T_898;
  wire [2:0] T_899;
  wire [8:0] T_900;
  wire [11:0] GEN_32;
  wire [11:0] T_901;
  reg [3:0] GEN_1;
  reg [31:0] GEN_41;
  assign io_req_ready = T_895;
  assign io_meta_read_valid = fire;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_1;
  assign io_meta_read_bits_tag = T_898;
  assign io_data_req_valid = fire;
  assign io_data_req_bits_way_en = req_way_en;
  assign io_data_req_bits_addr = T_901;
  assign io_release_valid = GEN_18;
  assign io_release_bits_addr_beat = beat_cnt;
  assign io_release_bits_addr_block = req_addr_block;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign io_release_bits_voluntary = req_voluntary;
  assign io_release_bits_r_type = req_r_type;
  assign io_release_bits_data = io_data_resp;
  assign T_748 = io_release_ready & io_release_valid;
  assign GEN_29 = {{2'd0}, 1'h1};
  assign T_753 = beat_cnt + GEN_29;
  assign T_754 = T_753[2:0];
  assign GEN_0 = T_748 ? T_754 : beat_cnt;
  assign T_864 = io_data_req_ready & io_data_req_valid;
  assign T_865 = io_meta_read_ready & io_meta_read_valid;
  assign T_866 = T_864 & T_865;
  assign GEN_30 = {{3'd0}, 1'h1};
  assign T_869 = data_req_cnt + GEN_30;
  assign T_870 = T_869[3:0];
  assign GEN_2 = T_866 ? T_870 : data_req_cnt;
  assign T_872 = io_release_ready == 1'h0;
  assign T_879 = r1_data_req_fired ? 2'h2 : {{1'd0}, 1'h1};
  assign GEN_31 = {{2'd0}, T_879};
  assign T_880 = data_req_cnt - GEN_31;
  assign T_881 = T_880[3:0];
  assign GEN_3 = T_872 ? 1'h0 : T_866;
  assign GEN_4 = T_872 ? 1'h0 : r1_data_req_fired;
  assign GEN_5 = T_872 ? T_881 : GEN_2;
  assign T_885 = r1_data_req_fired == 1'h0;
  assign T_887 = data_req_cnt < 4'h8;
  assign T_890 = T_887 | T_872;
  assign GEN_9 = T_885 ? T_890 : active;
  assign GEN_11 = r2_data_req_fired ? GEN_3 : T_866;
  assign GEN_12 = r2_data_req_fired ? GEN_4 : r1_data_req_fired;
  assign GEN_13 = r2_data_req_fired ? GEN_5 : GEN_2;
  assign GEN_14 = r2_data_req_fired ? GEN_9 : active;
  assign GEN_15 = active ? GEN_11 : r1_data_req_fired;
  assign GEN_16 = active ? GEN_12 : r2_data_req_fired;
  assign GEN_17 = active ? GEN_13 : data_req_cnt;
  assign GEN_18 = active ? r2_data_req_fired : 1'h0;
  assign GEN_19 = active ? GEN_14 : active;
  assign T_891 = io_req_ready & io_req_valid;
  assign GEN_20 = T_891 ? 1'h1 : GEN_19;
  assign GEN_21 = T_891 ? {{3'd0}, 1'h0} : GEN_17;
  assign GEN_22 = T_891 ? io_req_bits_addr_beat : req_addr_beat;
  assign GEN_23 = T_891 ? io_req_bits_addr_block : req_addr_block;
  assign GEN_24 = T_891 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign GEN_25 = T_891 ? io_req_bits_voluntary : req_voluntary;
  assign GEN_26 = T_891 ? io_req_bits_r_type : req_r_type;
  assign GEN_27 = T_891 ? io_req_bits_data : req_data;
  assign GEN_28 = T_891 ? io_req_bits_way_en : req_way_en;
  assign T_895 = active == 1'h0;
  assign req_idx = req_addr_block[5:0];
  assign fire = active & T_887;
  assign T_898 = req_addr_block[25:6];
  assign T_899 = data_req_cnt[2:0];
  assign T_900 = {req_idx,T_899};
  assign GEN_32 = {{3'd0}, T_900};
  assign T_901 = GEN_32 << 3;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_6 = {1{$random}};
  active = GEN_6[0:0];
  GEN_7 = {1{$random}};
  r1_data_req_fired = GEN_7[0:0];
  GEN_8 = {1{$random}};
  r2_data_req_fired = GEN_8[0:0];
  GEN_10 = {1{$random}};
  data_req_cnt = GEN_10[3:0];
  GEN_33 = {1{$random}};
  beat_cnt = GEN_33[2:0];
  GEN_34 = {1{$random}};
  req_addr_beat = GEN_34[2:0];
  GEN_35 = {1{$random}};
  req_addr_block = GEN_35[25:0];
  GEN_36 = {1{$random}};
  req_client_xact_id = GEN_36[1:0];
  GEN_37 = {1{$random}};
  req_voluntary = GEN_37[0:0];
  GEN_38 = {1{$random}};
  req_r_type = GEN_38[2:0];
  GEN_39 = {2{$random}};
  req_data = GEN_39[63:0];
  GEN_40 = {1{$random}};
  req_way_en = GEN_40[3:0];
  GEN_41 = {1{$random}};
  GEN_1 = GEN_41[3:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      active <= 1'h0;
    end else begin
      if(T_891) begin
        active <= 1'h1;
      end else begin
        if(active) begin
          if(r2_data_req_fired) begin
            if(T_885) begin
              active <= T_890;
            end
          end
        end
      end
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else begin
      if(active) begin
        if(r2_data_req_fired) begin
          if(T_872) begin
            r1_data_req_fired <= 1'h0;
          end else begin
            r1_data_req_fired <= T_866;
          end
        end else begin
          r1_data_req_fired <= T_866;
        end
      end
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else begin
      if(active) begin
        if(r2_data_req_fired) begin
          if(T_872) begin
            r2_data_req_fired <= 1'h0;
          end else begin
            r2_data_req_fired <= r1_data_req_fired;
          end
        end else begin
          r2_data_req_fired <= r1_data_req_fired;
        end
      end
    end
    if(reset) begin
      data_req_cnt <= 4'h0;
    end else begin
      if(T_891) begin
        data_req_cnt <= {{3'd0}, 1'h0};
      end else begin
        if(active) begin
          if(r2_data_req_fired) begin
            if(T_872) begin
              data_req_cnt <= T_881;
            end else begin
              if(T_866) begin
                data_req_cnt <= T_870;
              end
            end
          end else begin
            if(T_866) begin
              data_req_cnt <= T_870;
            end
          end
        end
      end
    end
    if(reset) begin
      beat_cnt <= 3'h0;
    end else begin
      if(T_748) begin
        beat_cnt <= T_754;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_891) begin
        req_addr_beat <= io_req_bits_addr_beat;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_891) begin
        req_addr_block <= io_req_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_891) begin
        req_client_xact_id <= io_req_bits_client_xact_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_891) begin
        req_voluntary <= io_req_bits_voluntary;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_891) begin
        req_r_type <= io_req_bits_r_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_891) begin
        req_data <= io_req_bits_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_891) begin
        req_way_en <= io_req_bits_way_en;
      end
    end
  end
endmodule
module ProbeUnit(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [25:0] io_req_bits_addr_block,
  input  [1:0] io_req_bits_p_type,
  input  [1:0] io_req_bits_client_xact_id,
  input   io_rep_ready,
  output  io_rep_valid,
  output [2:0] io_rep_bits_addr_beat,
  output [25:0] io_rep_bits_addr_block,
  output [1:0] io_rep_bits_client_xact_id,
  output  io_rep_bits_voluntary,
  output [2:0] io_rep_bits_r_type,
  output [63:0] io_rep_bits_data,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  input  [3:0] io_way_en,
  input   io_mshr_rdy,
  input  [1:0] io_block_state_state
);
  reg [3:0] state;
  reg [31:0] GEN_17;
  reg [1:0] old_coh_state;
  reg [31:0] GEN_18;
  reg [3:0] way_en;
  reg [31:0] GEN_19;
  reg [25:0] req_addr_block;
  reg [31:0] GEN_20;
  reg [1:0] req_p_type;
  reg [31:0] GEN_21;
  reg [1:0] req_client_xact_id;
  reg [31:0] GEN_22;
  wire [3:0] GEN_16;
  wire  tag_matches;
  wire [1:0] miss_coh_state;
  wire [1:0] reply_coh_state;
  wire [1:0] T_1256_0;
  wire  T_1258;
  wire [2:0] T_1261;
  wire [1:0] T_1275_0;
  wire  T_1277;
  wire [2:0] T_1281;
  wire [1:0] T_1294_0;
  wire  T_1296;
  wire [2:0] T_1301;
  wire  T_1308;
  wire [2:0] T_1309;
  wire  T_1310;
  wire [2:0] T_1311;
  wire  T_1312;
  wire [2:0] T_1313;
  wire [2:0] reply_addr_beat;
  wire [25:0] reply_addr_block;
  wire [1:0] reply_client_xact_id;
  wire  reply_voluntary;
  wire [2:0] reply_r_type;
  wire [63:0] reply_data;
  wire  T_1374;
  wire  T_1375;
  wire  T_1377;
  wire [2:0] T_1383_0;
  wire [2:0] T_1383_1;
  wire [2:0] T_1383_2;
  wire  T_1385;
  wire  T_1386;
  wire  T_1387;
  wire  T_1390;
  wire  T_1391;
  wire  T_1393;
  wire  T_1394;
  wire  T_1395;
  wire  T_1397;
  wire  T_1398;
  wire [19:0] T_1399;
  wire  T_1400;
  wire [1:0] T_1405;
  wire [1:0] T_1407;
  wire [1:0] T_1433_state;
  wire  T_1458;
  wire  T_1459;
  wire [3:0] GEN_0;
  wire [25:0] GEN_1;
  wire [1:0] GEN_2;
  wire [1:0] GEN_3;
  wire  T_1460;
  wire [3:0] GEN_4;
  wire  T_1461;
  wire [3:0] GEN_5;
  wire  T_1462;
  wire  T_1464;
  wire [3:0] GEN_6;
  wire [3:0] GEN_7;
  wire [1:0] GEN_8;
  wire [3:0] GEN_9;
  wire  T_1465;
  wire [1:0] T_1471_0;
  wire  T_1473;
  wire  T_1476;
  wire [3:0] T_1477;
  wire [3:0] GEN_11;
  wire  T_1479;
  wire [3:0] T_1480;
  wire [3:0] GEN_12;
  wire  T_1481;
  wire [3:0] GEN_13;
  wire  T_1482;
  wire  T_1483;
  wire [3:0] GEN_14;
  wire  T_1484;
  wire [3:0] GEN_15;
  reg [3:0] GEN_10;
  reg [31:0] GEN_23;
  assign io_req_ready = T_1374;
  assign io_rep_valid = T_1375;
  assign io_rep_bits_addr_beat = reply_addr_beat;
  assign io_rep_bits_addr_block = reply_addr_block;
  assign io_rep_bits_client_xact_id = reply_client_xact_id;
  assign io_rep_bits_voluntary = reply_voluntary;
  assign io_rep_bits_r_type = reply_r_type;
  assign io_rep_bits_data = reply_data;
  assign io_meta_read_valid = T_1398;
  assign io_meta_read_bits_idx = req_addr_block[5:0];
  assign io_meta_read_bits_way_en = GEN_10;
  assign io_meta_read_bits_tag = T_1399;
  assign io_meta_write_valid = T_1400;
  assign io_meta_write_bits_idx = req_addr_block[5:0];
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_data_tag = T_1399;
  assign io_meta_write_bits_data_coh_state = T_1433_state;
  assign io_wb_req_valid = T_1458;
  assign io_wb_req_bits_addr_beat = reply_addr_beat;
  assign io_wb_req_bits_addr_block = reply_addr_block;
  assign io_wb_req_bits_client_xact_id = reply_client_xact_id;
  assign io_wb_req_bits_voluntary = reply_voluntary;
  assign io_wb_req_bits_r_type = reply_r_type;
  assign io_wb_req_bits_data = reply_data;
  assign io_wb_req_bits_way_en = way_en;
  assign GEN_16 = {{3'd0}, 1'h0};
  assign tag_matches = way_en != GEN_16;
  assign miss_coh_state = {{1'd0}, 1'h0};
  assign reply_coh_state = tag_matches ? old_coh_state : miss_coh_state;
  assign T_1256_0 = 2'h3;
  assign T_1258 = T_1256_0 == reply_coh_state;
  assign T_1261 = T_1258 ? 3'h0 : 3'h3;
  assign T_1275_0 = 2'h3;
  assign T_1277 = T_1275_0 == reply_coh_state;
  assign T_1281 = T_1277 ? 3'h1 : 3'h4;
  assign T_1294_0 = 2'h3;
  assign T_1296 = T_1294_0 == reply_coh_state;
  assign T_1301 = T_1296 ? 3'h2 : 3'h5;
  assign T_1308 = 2'h2 == req_p_type;
  assign T_1309 = T_1308 ? T_1301 : 3'h3;
  assign T_1310 = 2'h1 == req_p_type;
  assign T_1311 = T_1310 ? T_1281 : T_1309;
  assign T_1312 = 2'h0 == req_p_type;
  assign T_1313 = T_1312 ? T_1261 : T_1311;
  assign reply_addr_beat = {{2'd0}, 1'h0};
  assign reply_addr_block = req_addr_block;
  assign reply_client_xact_id = {{1'd0}, 1'h0};
  assign reply_voluntary = 1'h0;
  assign reply_r_type = T_1313;
  assign reply_data = {{63'd0}, 1'h0};
  assign T_1374 = state == 4'h0;
  assign T_1375 = state == 4'h5;
  assign T_1377 = io_rep_valid == 1'h0;
  assign T_1383_0 = 3'h0;
  assign T_1383_1 = 3'h1;
  assign T_1383_2 = 3'h2;
  assign T_1385 = T_1383_0 == io_rep_bits_r_type;
  assign T_1386 = T_1383_1 == io_rep_bits_r_type;
  assign T_1387 = T_1383_2 == io_rep_bits_r_type;
  assign T_1390 = T_1385 | T_1386;
  assign T_1391 = T_1390 | T_1387;
  assign T_1393 = T_1391 == 1'h0;
  assign T_1394 = T_1377 | T_1393;
  assign T_1395 = T_1394 | reset;
  assign T_1397 = T_1395 == 1'h0;
  assign T_1398 = state == 4'h1;
  assign T_1399 = req_addr_block[25:6];
  assign T_1400 = state == 4'h8;
  assign T_1405 = T_1310 ? 2'h1 : old_coh_state;
  assign T_1407 = T_1312 ? 2'h0 : T_1405;
  assign T_1433_state = T_1407;
  assign T_1458 = state == 4'h6;
  assign T_1459 = io_req_ready & io_req_valid;
  assign GEN_0 = T_1459 ? 4'h1 : state;
  assign GEN_1 = T_1459 ? io_req_bits_addr_block : req_addr_block;
  assign GEN_2 = T_1459 ? io_req_bits_p_type : req_p_type;
  assign GEN_3 = T_1459 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign T_1460 = io_meta_read_ready & io_meta_read_valid;
  assign GEN_4 = T_1460 ? 4'h2 : GEN_0;
  assign T_1461 = state == 4'h2;
  assign GEN_5 = T_1461 ? 4'h3 : GEN_4;
  assign T_1462 = state == 4'h3;
  assign T_1464 = io_mshr_rdy == 1'h0;
  assign GEN_6 = T_1464 ? 4'h1 : 4'h4;
  assign GEN_7 = T_1462 ? GEN_6 : GEN_5;
  assign GEN_8 = T_1462 ? io_block_state_state : old_coh_state;
  assign GEN_9 = T_1462 ? io_way_en : way_en;
  assign T_1465 = state == 4'h4;
  assign T_1471_0 = 2'h3;
  assign T_1473 = T_1471_0 == old_coh_state;
  assign T_1476 = tag_matches & T_1473;
  assign T_1477 = T_1476 ? 4'h6 : 4'h5;
  assign GEN_11 = T_1465 ? T_1477 : GEN_7;
  assign T_1479 = T_1375 & io_rep_ready;
  assign T_1480 = tag_matches ? 4'h8 : 4'h0;
  assign GEN_12 = T_1479 ? T_1480 : GEN_11;
  assign T_1481 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_13 = T_1481 ? 4'h7 : GEN_12;
  assign T_1482 = state == 4'h7;
  assign T_1483 = T_1482 & io_wb_req_ready;
  assign GEN_14 = T_1483 ? 4'h8 : GEN_13;
  assign T_1484 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_15 = T_1484 ? 4'h0 : GEN_14;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_17 = {1{$random}};
  state = GEN_17[3:0];
  GEN_18 = {1{$random}};
  old_coh_state = GEN_18[1:0];
  GEN_19 = {1{$random}};
  way_en = GEN_19[3:0];
  GEN_20 = {1{$random}};
  req_addr_block = GEN_20[25:0];
  GEN_21 = {1{$random}};
  req_p_type = GEN_21[1:0];
  GEN_22 = {1{$random}};
  req_client_xact_id = GEN_22[1:0];
  GEN_23 = {1{$random}};
  GEN_10 = GEN_23[3:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_1484) begin
        state <= 4'h0;
      end else begin
        if(T_1483) begin
          state <= 4'h8;
        end else begin
          if(T_1481) begin
            state <= 4'h7;
          end else begin
            if(T_1479) begin
              if(tag_matches) begin
                state <= 4'h8;
              end else begin
                state <= 4'h0;
              end
            end else begin
              if(T_1465) begin
                if(T_1476) begin
                  state <= 4'h6;
                end else begin
                  state <= 4'h5;
                end
              end else begin
                if(T_1462) begin
                  if(T_1464) begin
                    state <= 4'h1;
                  end else begin
                    state <= 4'h4;
                  end
                end else begin
                  if(T_1461) begin
                    state <= 4'h3;
                  end else begin
                    if(T_1460) begin
                      state <= 4'h2;
                    end else begin
                      if(T_1459) begin
                        state <= 4'h1;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        old_coh_state <= io_block_state_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        way_en <= io_way_en;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1459) begin
        req_addr_block <= io_req_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1459) begin
        req_p_type <= io_req_bits_p_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1459) begin
        req_client_xact_id <= io_req_bits_client_xact_id;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1397) begin
          $fwrite(32'h80000002,"Assertion failed: ProbeUnit should not send releases with data\n    at nbdcache.scala:673 assert(!io.rep.valid || !io.rep.bits.hasData(),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1397) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1397) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Arbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  input  [19:0] io_in_0_bits_tag,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  input  [19:0] io_in_1_bits_tag,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [19:0] io_out_bits_tag,
  output  io_chosen
);
  wire  GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [19:0] GEN_3;
  wire  T_630;
  wire  T_632;
  wire  T_634;
  wire  T_635;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_632;
  assign io_out_valid = T_635;
  assign io_out_bits_idx = GEN_1;
  assign io_out_bits_way_en = GEN_2;
  assign io_out_bits_tag = GEN_3;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_idx : io_in_1_bits_idx;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag;
  assign T_630 = io_in_0_valid == 1'h0;
  assign T_632 = T_630 & io_out_ready;
  assign T_634 = T_630 == 1'h0;
  assign T_635 = T_634 | io_in_1_valid;
endmodule
module Arbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  input  [19:0] io_in_0_bits_data_tag,
  input  [1:0] io_in_0_bits_data_coh_state,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  input  [19:0] io_in_1_bits_data_tag,
  input  [1:0] io_in_1_bits_data_coh_state,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [19:0] io_out_bits_data_tag,
  output [1:0] io_out_bits_data_coh_state,
  output  io_chosen
);
  wire  GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [19:0] GEN_3;
  wire [1:0] GEN_4;
  wire  T_2720;
  wire  T_2722;
  wire  T_2724;
  wire  T_2725;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2722;
  assign io_out_valid = T_2725;
  assign io_out_bits_idx = GEN_1;
  assign io_out_bits_way_en = GEN_2;
  assign io_out_bits_data_tag = GEN_3;
  assign io_out_bits_data_coh_state = GEN_4;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_idx : io_in_1_bits_idx;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_data_coh_state : io_in_1_bits_data_coh_state;
  assign T_2720 = io_in_0_valid == 1'h0;
  assign T_2722 = T_2720 & io_out_ready;
  assign T_2724 = T_2720 == 1'h0;
  assign T_2725 = T_2724 | io_in_1_valid;
endmodule
module LockingArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [11:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [11:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_addr_beat,
  input   io_in_2_bits_is_builtin_type,
  input  [2:0] io_in_2_bits_a_type,
  input  [11:0] io_in_2_bits_union,
  input  [63:0] io_in_2_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [11:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire [1:0] GEN_29;
  wire  GEN_8;
  wire  GEN_9;
  wire [25:0] GEN_1;
  wire [25:0] GEN_10;
  wire [25:0] GEN_11;
  wire [1:0] GEN_2;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [2:0] GEN_3;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_4;
  wire  GEN_16;
  wire  GEN_17;
  wire [2:0] GEN_5;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [11:0] GEN_6;
  wire [11:0] GEN_20;
  wire [11:0] GEN_21;
  wire [63:0] GEN_7;
  wire [63:0] GEN_22;
  wire [63:0] GEN_23;
  reg [2:0] T_972;
  reg [31:0] GEN_30;
  reg [1:0] T_974;
  reg [31:0] GEN_31;
  wire [2:0] GEN_37;
  wire  T_976;
  wire [2:0] T_985_0;
  wire  T_987;
  wire  T_990;
  wire  T_991;
  wire  T_992;
  wire [2:0] GEN_38;
  wire [3:0] T_996;
  wire [2:0] T_997;
  wire [1:0] GEN_24;
  wire [2:0] GEN_25;
  wire [1:0] GEN_26;
  wire  T_999;
  wire  T_1001;
  wire  T_1003;
  wire [1:0] GEN_39;
  wire  T_1005;
  wire  T_1006;
  wire  T_1007;
  wire  T_1009;
  wire  T_1010;
  wire  T_1011;
  wire  T_1013;
  wire  T_1014;
  wire  T_1015;
  wire [1:0] GEN_27;
  wire [1:0] GEN_28;
  assign io_in_0_ready = T_1007;
  assign io_in_1_ready = T_1011;
  assign io_in_2_ready = T_1015;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_addr_beat = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_a_type = GEN_5;
  assign io_out_bits_union = GEN_6;
  assign io_out_bits_data = GEN_7;
  assign io_chosen = GEN_26;
  assign choice = GEN_28;
  assign GEN_0 = GEN_9;
  assign GEN_29 = {{1'd0}, 1'h1};
  assign GEN_8 = GEN_29 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_9 = 2'h2 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_1 = GEN_11;
  assign GEN_10 = GEN_29 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_10;
  assign GEN_2 = GEN_13;
  assign GEN_12 = GEN_29 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_12;
  assign GEN_3 = GEN_15;
  assign GEN_14 = GEN_29 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_14;
  assign GEN_4 = GEN_17;
  assign GEN_16 = GEN_29 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_16;
  assign GEN_5 = GEN_19;
  assign GEN_18 = GEN_29 == io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_a_type : GEN_18;
  assign GEN_6 = GEN_21;
  assign GEN_20 = GEN_29 == io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_union : GEN_20;
  assign GEN_7 = GEN_23;
  assign GEN_22 = GEN_29 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_22;
  assign GEN_37 = {{2'd0}, 1'h0};
  assign T_976 = T_972 != GEN_37;
  assign T_985_0 = 3'h3;
  assign T_987 = T_985_0 == io_out_bits_a_type;
  assign T_990 = io_out_bits_is_builtin_type & T_987;
  assign T_991 = io_out_ready & io_out_valid;
  assign T_992 = T_991 & T_990;
  assign GEN_38 = {{2'd0}, 1'h1};
  assign T_996 = T_972 + GEN_38;
  assign T_997 = T_996[2:0];
  assign GEN_24 = T_992 ? io_chosen : T_974;
  assign GEN_25 = T_992 ? T_997 : T_972;
  assign GEN_26 = T_976 ? T_974 : choice;
  assign T_999 = io_in_0_valid | io_in_1_valid;
  assign T_1001 = io_in_0_valid == 1'h0;
  assign T_1003 = T_999 == 1'h0;
  assign GEN_39 = {{1'd0}, 1'h0};
  assign T_1005 = T_974 == GEN_39;
  assign T_1006 = T_976 ? T_1005 : 1'h1;
  assign T_1007 = T_1006 & io_out_ready;
  assign T_1009 = T_974 == GEN_29;
  assign T_1010 = T_976 ? T_1009 : T_1001;
  assign T_1011 = T_1010 & io_out_ready;
  assign T_1013 = T_974 == 2'h2;
  assign T_1014 = T_976 ? T_1013 : T_1003;
  assign T_1015 = T_1014 & io_out_ready;
  assign GEN_27 = io_in_1_valid ? {{1'd0}, 1'h1} : 2'h2;
  assign GEN_28 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_27;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_30 = {1{$random}};
  T_972 = GEN_30[2:0];
  GEN_31 = {1{$random}};
  T_974 = GEN_31[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_972 <= 3'h0;
    end else begin
      if(T_992) begin
        T_972 <= T_997;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_992) begin
        T_974 <= io_chosen;
      end
    end
  end
endmodule
module Arbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_manager_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_manager_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_manager_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_manager_id,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [2:0] GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [2:0] GEN_4;
  wire  GEN_5;
  wire  T_716;
  wire  T_718;
  wire  T_720;
  wire  T_722;
  wire  T_723;
  wire  T_725;
  wire  T_726;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_722;
  assign io_in_2_ready = T_723;
  assign io_out_valid = T_726;
  assign io_out_bits_manager_xact_id = GEN_4;
  assign io_out_bits_manager_id = GEN_5;
  assign io_chosen = GEN_3;
  assign GEN_0 = io_in_1_valid ? {{1'd0}, 1'h1} : 2'h2;
  assign GEN_1 = io_in_1_valid ? io_in_1_bits_manager_xact_id : io_in_2_bits_manager_xact_id;
  assign GEN_2 = io_in_1_valid ? io_in_1_bits_manager_id : io_in_2_bits_manager_id;
  assign GEN_3 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_0;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_manager_xact_id : GEN_1;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_manager_id : GEN_2;
  assign T_716 = io_in_0_valid | io_in_1_valid;
  assign T_718 = io_in_0_valid == 1'h0;
  assign T_720 = T_716 == 1'h0;
  assign T_722 = T_718 & io_out_ready;
  assign T_723 = T_720 & io_out_ready;
  assign T_725 = T_720 == 1'h0;
  assign T_726 = T_725 | io_in_2_valid;
endmodule
module Arbiter_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  input  [3:0] io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  input  [3:0] io_in_1_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output [3:0] io_out_bits_way_en,
  output  io_chosen
);
  wire  GEN_0;
  wire [2:0] GEN_1;
  wire [25:0] GEN_2;
  wire [1:0] GEN_3;
  wire  GEN_4;
  wire [2:0] GEN_5;
  wire [63:0] GEN_6;
  wire [3:0] GEN_7;
  wire  T_1224;
  wire  T_1226;
  wire  T_1228;
  wire  T_1229;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1226;
  assign io_out_valid = T_1229;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_addr_block = GEN_2;
  assign io_out_bits_client_xact_id = GEN_3;
  assign io_out_bits_voluntary = GEN_4;
  assign io_out_bits_r_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_way_en = GEN_7;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr_beat : io_in_1_bits_addr_beat;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_addr_block : io_in_1_bits_addr_block;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_client_xact_id : io_in_1_bits_client_xact_id;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_voluntary : io_in_1_bits_voluntary;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_r_type : io_in_1_bits_r_type;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign T_1224 = io_in_0_valid == 1'h0;
  assign T_1226 = T_1224 & io_out_ready;
  assign T_1228 = T_1224 == 1'h0;
  assign T_1229 = T_1228 | io_in_1_valid;
endmodule
module Arbiter_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [8:0] io_in_0_bits_tag,
  input  [4:0] io_in_0_bits_cmd,
  input  [2:0] io_in_0_bits_typ,
  input   io_in_0_bits_phys,
  input  [4:0] io_in_0_bits_sdq_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [39:0] io_in_1_bits_addr,
  input  [8:0] io_in_1_bits_tag,
  input  [4:0] io_in_1_bits_cmd,
  input  [2:0] io_in_1_bits_typ,
  input   io_in_1_bits_phys,
  input  [4:0] io_in_1_bits_sdq_id,
  input   io_out_ready,
  output  io_out_valid,
  output [39:0] io_out_bits_addr,
  output [8:0] io_out_bits_tag,
  output [4:0] io_out_bits_cmd,
  output [2:0] io_out_bits_typ,
  output  io_out_bits_phys,
  output [4:0] io_out_bits_sdq_id,
  output  io_chosen
);
  wire  GEN_0;
  wire [39:0] GEN_1;
  wire [8:0] GEN_2;
  wire [4:0] GEN_3;
  wire [2:0] GEN_4;
  wire  GEN_5;
  wire [4:0] GEN_6;
  wire  T_1708;
  wire  T_1710;
  wire  T_1712;
  wire  T_1713;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1710;
  assign io_out_valid = T_1713;
  assign io_out_bits_addr = GEN_1;
  assign io_out_bits_tag = GEN_2;
  assign io_out_bits_cmd = GEN_3;
  assign io_out_bits_typ = GEN_4;
  assign io_out_bits_phys = GEN_5;
  assign io_out_bits_sdq_id = GEN_6;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_cmd : io_in_1_bits_cmd;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_typ : io_in_1_bits_typ;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_phys : io_in_1_bits_phys;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_sdq_id : io_in_1_bits_sdq_id;
  assign T_1708 = io_in_0_valid == 1'h0;
  assign T_1710 = T_1708 & io_out_ready;
  assign T_1712 = T_1708 == 1'h0;
  assign T_1713 = T_1712 | io_in_1_valid;
endmodule
module Arbiter_5(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input   io_in_1_bits,
  input   io_out_ready,
  output  io_out_valid,
  output  io_out_bits,
  output  io_chosen
);
  wire  GEN_0;
  wire  GEN_1;
  wire  T_58;
  wire  T_60;
  wire  T_62;
  wire  T_63;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_60;
  assign io_out_valid = T_63;
  assign io_out_bits = GEN_1;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits : io_in_1_bits;
  assign T_58 = io_in_0_valid == 1'h0;
  assign T_60 = T_58 & io_out_ready;
  assign T_62 = T_58 == 1'h0;
  assign T_63 = T_62 | io_in_1_valid;
endmodule
module Queue_1(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [39:0] io_enq_bits_addr,
  input  [8:0] io_enq_bits_tag,
  input  [4:0] io_enq_bits_cmd,
  input  [2:0] io_enq_bits_typ,
  input   io_enq_bits_phys,
  input  [4:0] io_enq_bits_sdq_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [39:0] io_deq_bits_addr,
  output [8:0] io_deq_bits_tag,
  output [4:0] io_deq_bits_cmd,
  output [2:0] io_deq_bits_typ,
  output  io_deq_bits_phys,
  output [4:0] io_deq_bits_sdq_id,
  output [4:0] io_count
);
  reg [39:0] ram_addr [0:15];
  reg [63:0] GEN_0;
  wire [39:0] ram_addr_T_794_data;
  wire [3:0] ram_addr_T_794_addr;
  wire  ram_addr_T_794_en;
  wire [39:0] ram_addr_T_703_data;
  wire [3:0] ram_addr_T_703_addr;
  wire  ram_addr_T_703_mask;
  wire  ram_addr_T_703_en;
  reg [8:0] ram_tag [0:15];
  reg [31:0] GEN_1;
  wire [8:0] ram_tag_T_794_data;
  wire [3:0] ram_tag_T_794_addr;
  wire  ram_tag_T_794_en;
  wire [8:0] ram_tag_T_703_data;
  wire [3:0] ram_tag_T_703_addr;
  wire  ram_tag_T_703_mask;
  wire  ram_tag_T_703_en;
  reg [4:0] ram_cmd [0:15];
  reg [31:0] GEN_2;
  wire [4:0] ram_cmd_T_794_data;
  wire [3:0] ram_cmd_T_794_addr;
  wire  ram_cmd_T_794_en;
  wire [4:0] ram_cmd_T_703_data;
  wire [3:0] ram_cmd_T_703_addr;
  wire  ram_cmd_T_703_mask;
  wire  ram_cmd_T_703_en;
  reg [2:0] ram_typ [0:15];
  reg [31:0] GEN_3;
  wire [2:0] ram_typ_T_794_data;
  wire [3:0] ram_typ_T_794_addr;
  wire  ram_typ_T_794_en;
  wire [2:0] ram_typ_T_703_data;
  wire [3:0] ram_typ_T_703_addr;
  wire  ram_typ_T_703_mask;
  wire  ram_typ_T_703_en;
  reg  ram_phys [0:15];
  reg [31:0] GEN_4;
  wire  ram_phys_T_794_data;
  wire [3:0] ram_phys_T_794_addr;
  wire  ram_phys_T_794_en;
  wire  ram_phys_T_703_data;
  wire [3:0] ram_phys_T_703_addr;
  wire  ram_phys_T_703_mask;
  wire  ram_phys_T_703_en;
  reg [4:0] ram_sdq_id [0:15];
  reg [31:0] GEN_5;
  wire [4:0] ram_sdq_id_T_794_data;
  wire [3:0] ram_sdq_id_T_794_addr;
  wire  ram_sdq_id_T_794_en;
  wire [4:0] ram_sdq_id_T_703_data;
  wire [3:0] ram_sdq_id_T_703_addr;
  wire  ram_sdq_id_T_703_mask;
  wire  ram_sdq_id_T_703_en;
  reg [3:0] T_695;
  reg [31:0] GEN_6;
  reg [3:0] T_697;
  reg [31:0] GEN_7;
  reg  maybe_full;
  reg [31:0] GEN_8;
  wire  ptr_match;
  wire  T_700;
  wire  empty;
  wire  full;
  wire  T_701;
  wire  do_enq;
  wire  T_702;
  wire  do_deq;
  wire [3:0] GEN_18;
  wire [4:0] T_782;
  wire [3:0] T_783;
  wire [3:0] GEN_15;
  wire [4:0] T_787;
  wire [3:0] T_788;
  wire [3:0] GEN_16;
  wire  T_789;
  wire  GEN_17;
  wire  T_791;
  wire  T_793;
  wire [4:0] T_870;
  wire [3:0] ptr_diff;
  wire  T_871;
  wire [4:0] T_872;
  assign io_enq_ready = T_793;
  assign io_deq_valid = T_791;
  assign io_deq_bits_addr = ram_addr_T_794_data;
  assign io_deq_bits_tag = ram_tag_T_794_data;
  assign io_deq_bits_cmd = ram_cmd_T_794_data;
  assign io_deq_bits_typ = ram_typ_T_794_data;
  assign io_deq_bits_phys = ram_phys_T_794_data;
  assign io_deq_bits_sdq_id = ram_sdq_id_T_794_data;
  assign io_count = T_872;
  assign ram_addr_T_794_addr = T_697;
  assign ram_addr_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_T_794_data = ram_addr[ram_addr_T_794_addr];
  `else
  assign ram_addr_T_794_data = ram_addr_T_794_addr >= 5'h10 ? $random : ram_addr[ram_addr_T_794_addr];
  `endif
  assign ram_addr_T_703_data = io_enq_bits_addr;
  assign ram_addr_T_703_addr = T_695;
  assign ram_addr_T_703_mask = do_enq;
  assign ram_addr_T_703_en = do_enq;
  assign ram_tag_T_794_addr = T_697;
  assign ram_tag_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_tag_T_794_data = ram_tag[ram_tag_T_794_addr];
  `else
  assign ram_tag_T_794_data = ram_tag_T_794_addr >= 5'h10 ? $random : ram_tag[ram_tag_T_794_addr];
  `endif
  assign ram_tag_T_703_data = io_enq_bits_tag;
  assign ram_tag_T_703_addr = T_695;
  assign ram_tag_T_703_mask = do_enq;
  assign ram_tag_T_703_en = do_enq;
  assign ram_cmd_T_794_addr = T_697;
  assign ram_cmd_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_cmd_T_794_data = ram_cmd[ram_cmd_T_794_addr];
  `else
  assign ram_cmd_T_794_data = ram_cmd_T_794_addr >= 5'h10 ? $random : ram_cmd[ram_cmd_T_794_addr];
  `endif
  assign ram_cmd_T_703_data = io_enq_bits_cmd;
  assign ram_cmd_T_703_addr = T_695;
  assign ram_cmd_T_703_mask = do_enq;
  assign ram_cmd_T_703_en = do_enq;
  assign ram_typ_T_794_addr = T_697;
  assign ram_typ_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_typ_T_794_data = ram_typ[ram_typ_T_794_addr];
  `else
  assign ram_typ_T_794_data = ram_typ_T_794_addr >= 5'h10 ? $random : ram_typ[ram_typ_T_794_addr];
  `endif
  assign ram_typ_T_703_data = io_enq_bits_typ;
  assign ram_typ_T_703_addr = T_695;
  assign ram_typ_T_703_mask = do_enq;
  assign ram_typ_T_703_en = do_enq;
  assign ram_phys_T_794_addr = T_697;
  assign ram_phys_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_phys_T_794_data = ram_phys[ram_phys_T_794_addr];
  `else
  assign ram_phys_T_794_data = ram_phys_T_794_addr >= 5'h10 ? $random : ram_phys[ram_phys_T_794_addr];
  `endif
  assign ram_phys_T_703_data = io_enq_bits_phys;
  assign ram_phys_T_703_addr = T_695;
  assign ram_phys_T_703_mask = do_enq;
  assign ram_phys_T_703_en = do_enq;
  assign ram_sdq_id_T_794_addr = T_697;
  assign ram_sdq_id_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_sdq_id_T_794_data = ram_sdq_id[ram_sdq_id_T_794_addr];
  `else
  assign ram_sdq_id_T_794_data = ram_sdq_id_T_794_addr >= 5'h10 ? $random : ram_sdq_id[ram_sdq_id_T_794_addr];
  `endif
  assign ram_sdq_id_T_703_data = io_enq_bits_sdq_id;
  assign ram_sdq_id_T_703_addr = T_695;
  assign ram_sdq_id_T_703_mask = do_enq;
  assign ram_sdq_id_T_703_en = do_enq;
  assign ptr_match = T_695 == T_697;
  assign T_700 = maybe_full == 1'h0;
  assign empty = ptr_match & T_700;
  assign full = ptr_match & maybe_full;
  assign T_701 = io_enq_ready & io_enq_valid;
  assign do_enq = T_701;
  assign T_702 = io_deq_ready & io_deq_valid;
  assign do_deq = T_702;
  assign GEN_18 = {{3'd0}, 1'h1};
  assign T_782 = T_695 + GEN_18;
  assign T_783 = T_782[3:0];
  assign GEN_15 = do_enq ? T_783 : T_695;
  assign T_787 = T_697 + GEN_18;
  assign T_788 = T_787[3:0];
  assign GEN_16 = do_deq ? T_788 : T_697;
  assign T_789 = do_enq != do_deq;
  assign GEN_17 = T_789 ? do_enq : maybe_full;
  assign T_791 = empty == 1'h0;
  assign T_793 = full == 1'h0;
  assign T_870 = T_695 - T_697;
  assign ptr_diff = T_870[3:0];
  assign T_871 = maybe_full & ptr_match;
  assign T_872 = {T_871,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {2{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_addr[initvar] = GEN_0[39:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_tag[initvar] = GEN_1[8:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_cmd[initvar] = GEN_2[4:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_typ[initvar] = GEN_3[2:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_phys[initvar] = GEN_4[0:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_sdq_id[initvar] = GEN_5[4:0];
  GEN_6 = {1{$random}};
  T_695 = GEN_6[3:0];
  GEN_7 = {1{$random}};
  T_697 = GEN_7[3:0];
  GEN_8 = {1{$random}};
  maybe_full = GEN_8[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_T_703_en & ram_addr_T_703_mask) begin
      ram_addr[ram_addr_T_703_addr] <= ram_addr_T_703_data;
    end
    if(ram_tag_T_703_en & ram_tag_T_703_mask) begin
      ram_tag[ram_tag_T_703_addr] <= ram_tag_T_703_data;
    end
    if(ram_cmd_T_703_en & ram_cmd_T_703_mask) begin
      ram_cmd[ram_cmd_T_703_addr] <= ram_cmd_T_703_data;
    end
    if(ram_typ_T_703_en & ram_typ_T_703_mask) begin
      ram_typ[ram_typ_T_703_addr] <= ram_typ_T_703_data;
    end
    if(ram_phys_T_703_en & ram_phys_T_703_mask) begin
      ram_phys[ram_phys_T_703_addr] <= ram_phys_T_703_data;
    end
    if(ram_sdq_id_T_703_en & ram_sdq_id_T_703_mask) begin
      ram_sdq_id[ram_sdq_id_T_703_addr] <= ram_sdq_id_T_703_data;
    end
    if(reset) begin
      T_695 <= 4'h0;
    end else begin
      if(do_enq) begin
        T_695 <= T_783;
      end
    end
    if(reset) begin
      T_697 <= 4'h0;
    end else begin
      if(do_deq) begin
        T_697 <= T_788;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_789) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module FinishQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output  io_count
);
  reg [2:0] T_244_manager_xact_id [0:0];
  reg [31:0] GEN_0;
  wire [2:0] T_244_manager_xact_id_T_291_data;
  wire  T_244_manager_xact_id_T_291_addr;
  wire  T_244_manager_xact_id_T_291_en;
  wire [2:0] T_244_manager_xact_id_T_258_data;
  wire  T_244_manager_xact_id_T_258_addr;
  wire  T_244_manager_xact_id_T_258_mask;
  wire  T_244_manager_xact_id_T_258_en;
  reg  T_244_manager_id [0:0];
  reg [31:0] GEN_1;
  wire  T_244_manager_id_T_291_data;
  wire  T_244_manager_id_T_291_addr;
  wire  T_244_manager_id_T_291_en;
  wire  T_244_manager_id_T_258_data;
  wire  T_244_manager_id_T_258_addr;
  wire  T_244_manager_id_T_258_mask;
  wire  T_244_manager_id_T_258_en;
  reg  T_248;
  reg [31:0] GEN_2;
  wire  T_251;
  wire  T_254;
  wire  T_255;
  wire  T_256;
  wire  T_257;
  wire  T_286;
  wire  GEN_7;
  wire  T_288;
  wire [1:0] T_317;
  wire  T_318;
  wire [1:0] T_320;
  assign io_enq_ready = T_251;
  assign io_deq_valid = T_288;
  assign io_deq_bits_manager_xact_id = T_244_manager_xact_id_T_291_data;
  assign io_deq_bits_manager_id = T_244_manager_id_T_291_data;
  assign io_count = T_320[0];
  assign T_244_manager_xact_id_T_291_addr = 1'h0;
  assign T_244_manager_xact_id_T_291_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_244_manager_xact_id_T_291_data = T_244_manager_xact_id[T_244_manager_xact_id_T_291_addr];
  `else
  assign T_244_manager_xact_id_T_291_data = T_244_manager_xact_id_T_291_addr >= 1'h1 ? $random : T_244_manager_xact_id[T_244_manager_xact_id_T_291_addr];
  `endif
  assign T_244_manager_xact_id_T_258_data = io_enq_bits_manager_xact_id;
  assign T_244_manager_xact_id_T_258_addr = 1'h0;
  assign T_244_manager_xact_id_T_258_mask = T_255;
  assign T_244_manager_xact_id_T_258_en = T_255;
  assign T_244_manager_id_T_291_addr = 1'h0;
  assign T_244_manager_id_T_291_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_244_manager_id_T_291_data = T_244_manager_id[T_244_manager_id_T_291_addr];
  `else
  assign T_244_manager_id_T_291_data = T_244_manager_id_T_291_addr >= 1'h1 ? $random : T_244_manager_id[T_244_manager_id_T_291_addr];
  `endif
  assign T_244_manager_id_T_258_data = io_enq_bits_manager_id;
  assign T_244_manager_id_T_258_addr = 1'h0;
  assign T_244_manager_id_T_258_mask = T_255;
  assign T_244_manager_id_T_258_en = T_255;
  assign T_251 = T_248 == 1'h0;
  assign T_254 = io_enq_ready & io_enq_valid;
  assign T_255 = T_254;
  assign T_256 = io_deq_ready & io_deq_valid;
  assign T_257 = T_256;
  assign T_286 = T_255 != T_257;
  assign GEN_7 = T_286 ? T_255 : T_248;
  assign T_288 = T_251 == 1'h0;
  assign T_317 = 1'h0 - 1'h0;
  assign T_318 = T_317[0:0];
  assign T_320 = {T_248,T_318};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    T_244_manager_xact_id[initvar] = GEN_0[2:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    T_244_manager_id[initvar] = GEN_1[0:0];
  GEN_2 = {1{$random}};
  T_248 = GEN_2[0:0];
  end
`endif
  always @(posedge clk) begin
    if(T_244_manager_xact_id_T_258_en & T_244_manager_xact_id_T_258_mask) begin
      T_244_manager_xact_id[T_244_manager_xact_id_T_258_addr] <= T_244_manager_xact_id_T_258_data;
    end
    if(T_244_manager_id_T_258_en & T_244_manager_id_T_258_mask) begin
      T_244_manager_id[T_244_manager_id_T_258_addr] <= T_244_manager_id_T_258_data;
    end
    if(reset) begin
      T_248 <= 1'h0;
    end else begin
      if(T_286) begin
        T_248 <= T_255;
      end
    end
  end
endmodule
module MSHR(
  input   clk,
  input   reset,
  input   io_req_pri_val,
  output  io_req_pri_rdy,
  input   io_req_sec_val,
  output  io_req_sec_rdy,
  input  [39:0] io_req_bits_addr,
  input  [8:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [4:0] io_req_bits_sdq_id,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  output  io_idx_match,
  output [19:0] io_tag,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [11:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [8:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [4:0] io_replay_bits_sdq_id,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy
);
  reg [3:0] state;
  reg [31:0] GEN_16;
  wire [1:0] T_1875_state;
  reg [1:0] new_coh_state_state;
  reg [31:0] GEN_17;
  reg [39:0] req_addr;
  reg [63:0] GEN_18;
  reg [8:0] req_tag;
  reg [31:0] GEN_19;
  reg [4:0] req_cmd;
  reg [31:0] GEN_22;
  reg [2:0] req_typ;
  reg [31:0] GEN_34;
  reg  req_phys;
  reg [31:0] GEN_35;
  reg [4:0] req_sdq_id;
  reg [31:0] GEN_36;
  reg  req_tag_match;
  reg [31:0] GEN_37;
  reg [19:0] req_old_meta_tag;
  reg [31:0] GEN_38;
  reg [1:0] req_old_meta_coh_state;
  reg [31:0] GEN_41;
  reg [3:0] req_way_en;
  reg [31:0] GEN_57;
  wire [5:0] req_idx;
  wire [5:0] T_2271;
  wire  idx_match;
  wire  T_2272;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2278;
  wire  T_2279;
  wire  T_2280;
  wire  T_2281;
  wire  T_2282;
  wire  T_2283;
  wire  T_2284;
  wire  T_2285;
  wire  T_2286;
  wire  T_2287;
  wire  T_2288;
  wire  T_2289;
  wire  T_2290;
  wire  T_2291;
  wire  T_2292;
  wire  T_2293;
  wire  T_2295;
  wire  cmd_requires_second_acquire;
  wire [3:0] states_before_refill_0;
  wire [3:0] states_before_refill_1;
  wire [3:0] states_before_refill_2;
  wire  T_2302;
  wire  T_2303;
  wire  T_2304;
  wire  T_2307;
  wire  T_2308;
  wire [3:0] T_2314_0;
  wire [3:0] T_2314_1;
  wire  T_2316;
  wire  T_2317;
  wire  T_2320;
  wire  T_2322;
  wire  T_2323;
  wire  T_2324;
  wire  sec_rdy;
  wire [2:0] T_2332_0;
  wire [3:0] GEN_46;
  wire  T_2334;
  wire [1:0] T_2342_0;
  wire [1:0] T_2342_1;
  wire [3:0] GEN_47;
  wire  T_2344;
  wire [3:0] GEN_48;
  wire  T_2345;
  wire  T_2348;
  wire  T_2349;
  wire  T_2350;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_58;
  wire  T_2353;
  wire [2:0] GEN_49;
  wire [3:0] T_2355;
  wire [2:0] T_2356;
  wire [2:0] GEN_0;
  wire  refill_count_done;
  wire  T_2358;
  wire  T_2359;
  wire  refill_done;
  wire  rpq_clk;
  wire  rpq_reset;
  wire  rpq_io_enq_ready;
  wire  rpq_io_enq_valid;
  wire [39:0] rpq_io_enq_bits_addr;
  wire [8:0] rpq_io_enq_bits_tag;
  wire [4:0] rpq_io_enq_bits_cmd;
  wire [2:0] rpq_io_enq_bits_typ;
  wire  rpq_io_enq_bits_phys;
  wire [4:0] rpq_io_enq_bits_sdq_id;
  wire  rpq_io_deq_ready;
  wire  rpq_io_deq_valid;
  wire [39:0] rpq_io_deq_bits_addr;
  wire [8:0] rpq_io_deq_bits_tag;
  wire [4:0] rpq_io_deq_bits_cmd;
  wire [2:0] rpq_io_deq_bits_typ;
  wire  rpq_io_deq_bits_phys;
  wire [4:0] rpq_io_deq_bits_sdq_id;
  wire [4:0] rpq_io_count;
  wire  T_2436;
  wire  T_2437;
  wire  T_2438;
  wire  T_2439;
  wire  T_2441;
  wire  T_2443;
  wire  T_2444;
  wire  T_2445;
  wire  T_2446;
  wire  T_2447;
  wire  T_2448;
  wire [1:0] T_2456;
  wire [3:0] GEN_50;
  wire  T_2457;
  wire [1:0] T_2458;
  wire [3:0] GEN_51;
  wire  T_2459;
  wire [1:0] T_2460;
  wire [3:0] GEN_52;
  wire  T_2461;
  wire [1:0] T_2462;
  wire [1:0] T_2463;
  wire [1:0] coh_on_grant_state;
  wire [1:0] T_2520;
  wire [1:0] coh_on_hit_state;
  wire  T_2572;
  wire  T_2573;
  wire [3:0] GEN_1;
  wire  T_2574;
  wire [3:0] GEN_2;
  wire  T_2575;
  wire  T_2576;
  wire [3:0] GEN_3;
  wire  T_2577;
  wire  T_2578;
  wire [3:0] GEN_4;
  wire [1:0] GEN_5;
  wire  T_2579;
  wire [3:0] GEN_6;
  wire  T_2580;
  wire  T_2581;
  wire [3:0] GEN_7;
  wire  T_2582;
  wire  T_2583;
  wire [3:0] GEN_8;
  wire  T_2584;
  wire [3:0] GEN_9;
  wire  T_2589;
  wire [4:0] GEN_10;
  wire [4:0] GEN_11;
  wire [1:0] T_2607_0;
  wire [1:0] T_2607_1;
  wire  T_2609;
  wire  T_2610;
  wire  T_2613;
  wire [1:0] T_2619_0;
  wire [1:0] T_2619_1;
  wire [1:0] T_2619_2;
  wire  T_2621;
  wire  T_2622;
  wire  T_2623;
  wire  T_2626;
  wire  T_2627;
  wire  T_2628;
  wire [3:0] GEN_12;
  wire [1:0] GEN_13;
  wire  T_2630;
  wire [3:0] GEN_14;
  wire [3:0] GEN_20;
  wire [1:0] GEN_21;
  wire  T_2632;
  wire [1:0] T_2638_0;
  wire  T_2640;
  wire [3:0] T_2643;
  wire [3:0] GEN_23;
  wire [39:0] GEN_24;
  wire [8:0] GEN_25;
  wire [4:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [4:0] GEN_29;
  wire  GEN_30;
  wire [19:0] GEN_31;
  wire [1:0] GEN_32;
  wire [3:0] GEN_33;
  wire [3:0] GEN_39;
  wire [1:0] GEN_40;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  wire  T_2671;
  wire  can_finish;
  wire [3:0] GEN_53;
  wire  T_2676;
  wire  T_2677;
  wire  T_2679;
  wire  T_2681;
  wire  T_2682;
  wire [2:0] T_2709_manager_xact_id;
  wire  T_2709_manager_id;
  wire  T_2735;
  wire  T_2736;
  wire  T_2737;
  wire  T_2738;
  wire [8:0] T_2739;
  wire [11:0] GEN_54;
  wire [11:0] T_2740;
  wire [27:0] T_2741;
  wire  T_2743;
  reg [1:0] meta_hazard;
  reg [31:0] GEN_59;
  wire [1:0] GEN_55;
  wire  T_2746;
  wire [1:0] GEN_56;
  wire [2:0] T_2748;
  wire [1:0] T_2749;
  wire [1:0] GEN_42;
  wire  T_2750;
  wire [1:0] GEN_43;
  wire  T_2753;
  wire  T_2762;
  wire  T_2764;
  wire  T_2765;
  wire  T_2766;
  wire  T_2769;
  wire [1:0] T_2776_0;
  wire [1:0] T_2776_1;
  wire [1:0] T_2817_state;
  wire [1:0] T_2842_state;
  wire  T_2867;
  wire [25:0] T_2869;
  wire [1:0] T_2878_0;
  wire  T_2880;
  wire [2:0] T_2883;
  wire [2:0] T_2922_addr_beat;
  wire [25:0] T_2922_addr_block;
  wire [1:0] T_2922_client_xact_id;
  wire  T_2922_voluntary;
  wire [2:0] T_2922_r_type;
  wire [63:0] T_2922_data;
  wire  T_2953;
  wire [25:0] T_2954;
  wire [5:0] T_2970;
  wire [25:0] T_3004_addr_block;
  wire [1:0] T_3004_client_xact_id;
  wire [2:0] T_3004_addr_beat;
  wire  T_3004_is_builtin_type;
  wire [2:0] T_3004_a_type;
  wire [11:0] T_3004_union;
  wire [63:0] T_3004_data;
  wire  T_3037;
  wire [5:0] T_3039;
  wire [31:0] T_3041;
  wire  T_3043;
  wire  GEN_44;
  wire [4:0] GEN_45;
  reg [3:0] GEN_15;
  reg [31:0] GEN_60;
  Queue_1 rpq (
    .clk(rpq_clk),
    .reset(rpq_reset),
    .io_enq_ready(rpq_io_enq_ready),
    .io_enq_valid(rpq_io_enq_valid),
    .io_enq_bits_addr(rpq_io_enq_bits_addr),
    .io_enq_bits_tag(rpq_io_enq_bits_tag),
    .io_enq_bits_cmd(rpq_io_enq_bits_cmd),
    .io_enq_bits_typ(rpq_io_enq_bits_typ),
    .io_enq_bits_phys(rpq_io_enq_bits_phys),
    .io_enq_bits_sdq_id(rpq_io_enq_bits_sdq_id),
    .io_deq_ready(rpq_io_deq_ready),
    .io_deq_valid(rpq_io_deq_valid),
    .io_deq_bits_addr(rpq_io_deq_bits_addr),
    .io_deq_bits_tag(rpq_io_deq_bits_tag),
    .io_deq_bits_cmd(rpq_io_deq_bits_cmd),
    .io_deq_bits_typ(rpq_io_deq_bits_typ),
    .io_deq_bits_phys(rpq_io_deq_bits_phys),
    .io_deq_bits_sdq_id(rpq_io_deq_bits_sdq_id),
    .io_count(rpq_io_count)
  );
  FinishQueue fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_pri_rdy = T_2447;
  assign io_req_sec_rdy = T_2743;
  assign io_idx_match = T_2738;
  assign io_tag = T_2741[19:0];
  assign io_mem_req_valid = T_2953;
  assign io_mem_req_bits_addr_block = T_3004_addr_block;
  assign io_mem_req_bits_client_xact_id = T_3004_client_xact_id;
  assign io_mem_req_bits_addr_beat = T_3004_addr_beat;
  assign io_mem_req_bits_is_builtin_type = T_3004_is_builtin_type;
  assign io_mem_req_bits_a_type = T_3004_a_type;
  assign io_mem_req_bits_union = T_3004_union;
  assign io_mem_req_bits_data = T_3004_data;
  assign io_refill_way_en = req_way_en;
  assign io_refill_addr = T_2740;
  assign io_meta_read_valid = T_2445;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_15;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_write_valid = T_2769;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_data_coh_state = T_2842_state;
  assign io_replay_valid = T_3037;
  assign io_replay_bits_addr = {{8'd0}, T_3041};
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_cmd = GEN_45;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_mem_finish_valid = T_2735;
  assign io_mem_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_wb_req_valid = T_2867;
  assign io_wb_req_bits_addr_beat = T_2922_addr_beat;
  assign io_wb_req_bits_addr_block = T_2922_addr_block;
  assign io_wb_req_bits_client_xact_id = T_2922_client_xact_id;
  assign io_wb_req_bits_voluntary = T_2922_voluntary;
  assign io_wb_req_bits_r_type = T_2922_r_type;
  assign io_wb_req_bits_data = T_2922_data;
  assign io_wb_req_bits_way_en = req_way_en;
  assign io_probe_rdy = T_2766;
  assign T_1875_state = {{1'd0}, 1'h0};
  assign req_idx = req_addr[11:6];
  assign T_2271 = io_req_bits_addr[11:6];
  assign idx_match = req_idx == T_2271;
  assign T_2272 = io_req_bits_cmd == 5'h1;
  assign T_2273 = io_req_bits_cmd == 5'h7;
  assign T_2274 = T_2272 | T_2273;
  assign T_2275 = io_req_bits_cmd[3];
  assign T_2276 = io_req_bits_cmd == 5'h4;
  assign T_2277 = T_2275 | T_2276;
  assign T_2278 = T_2274 | T_2277;
  assign T_2279 = io_req_bits_cmd == 5'h3;
  assign T_2280 = T_2278 | T_2279;
  assign T_2281 = io_req_bits_cmd == 5'h6;
  assign T_2282 = T_2280 | T_2281;
  assign T_2283 = req_cmd == 5'h1;
  assign T_2284 = req_cmd == 5'h7;
  assign T_2285 = T_2283 | T_2284;
  assign T_2286 = req_cmd[3];
  assign T_2287 = req_cmd == 5'h4;
  assign T_2288 = T_2286 | T_2287;
  assign T_2289 = T_2285 | T_2288;
  assign T_2290 = req_cmd == 5'h3;
  assign T_2291 = T_2289 | T_2290;
  assign T_2292 = req_cmd == 5'h6;
  assign T_2293 = T_2291 | T_2292;
  assign T_2295 = T_2293 == 1'h0;
  assign cmd_requires_second_acquire = T_2282 & T_2295;
  assign states_before_refill_0 = 4'h1;
  assign states_before_refill_1 = 4'h2;
  assign states_before_refill_2 = 4'h3;
  assign T_2302 = states_before_refill_0 == state;
  assign T_2303 = states_before_refill_1 == state;
  assign T_2304 = states_before_refill_2 == state;
  assign T_2307 = T_2302 | T_2303;
  assign T_2308 = T_2307 | T_2304;
  assign T_2314_0 = 4'h4;
  assign T_2314_1 = 4'h5;
  assign T_2316 = T_2314_0 == state;
  assign T_2317 = T_2314_1 == state;
  assign T_2320 = T_2316 | T_2317;
  assign T_2322 = cmd_requires_second_acquire == 1'h0;
  assign T_2323 = T_2320 & T_2322;
  assign T_2324 = T_2308 | T_2323;
  assign sec_rdy = idx_match & T_2324;
  assign T_2332_0 = 3'h5;
  assign GEN_46 = {{1'd0}, T_2332_0};
  assign T_2334 = GEN_46 == io_mem_grant_bits_g_type;
  assign T_2342_0 = 2'h0;
  assign T_2342_1 = 2'h1;
  assign GEN_47 = {{2'd0}, T_2342_0};
  assign T_2344 = GEN_47 == io_mem_grant_bits_g_type;
  assign GEN_48 = {{2'd0}, T_2342_1};
  assign T_2345 = GEN_48 == io_mem_grant_bits_g_type;
  assign T_2348 = T_2344 | T_2345;
  assign T_2349 = io_mem_grant_bits_is_builtin_type ? T_2334 : T_2348;
  assign T_2350 = io_mem_grant_valid & T_2349;
  assign T_2353 = refill_cnt == 3'h7;
  assign GEN_49 = {{2'd0}, 1'h1};
  assign T_2355 = refill_cnt + GEN_49;
  assign T_2356 = T_2355[2:0];
  assign GEN_0 = T_2350 ? T_2356 : refill_cnt;
  assign refill_count_done = T_2350 & T_2353;
  assign T_2358 = T_2349 == 1'h0;
  assign T_2359 = T_2358 | refill_count_done;
  assign refill_done = io_mem_grant_valid & T_2359;
  assign rpq_clk = clk;
  assign rpq_reset = reset;
  assign rpq_io_enq_valid = T_2444;
  assign rpq_io_enq_bits_addr = io_req_bits_addr;
  assign rpq_io_enq_bits_tag = io_req_bits_tag;
  assign rpq_io_enq_bits_cmd = io_req_bits_cmd;
  assign rpq_io_enq_bits_typ = io_req_bits_typ;
  assign rpq_io_enq_bits_phys = io_req_bits_phys;
  assign rpq_io_enq_bits_sdq_id = io_req_bits_sdq_id;
  assign rpq_io_deq_ready = GEN_44;
  assign T_2436 = io_req_pri_val & io_req_pri_rdy;
  assign T_2437 = io_req_sec_val & sec_rdy;
  assign T_2438 = T_2436 | T_2437;
  assign T_2439 = io_req_bits_cmd == 5'h2;
  assign T_2441 = T_2439 | T_2279;
  assign T_2443 = T_2441 == 1'h0;
  assign T_2444 = T_2438 & T_2443;
  assign T_2445 = state == 4'h8;
  assign T_2446 = io_replay_ready & T_2445;
  assign T_2447 = state == 4'h0;
  assign T_2448 = T_2446 | T_2447;
  assign T_2456 = T_2289 ? 2'h3 : 2'h2;
  assign GEN_50 = {{2'd0}, 2'h2};
  assign T_2457 = GEN_50 == io_mem_grant_bits_g_type;
  assign T_2458 = T_2457 ? 2'h3 : 2'h0;
  assign GEN_51 = {{2'd0}, 2'h1};
  assign T_2459 = GEN_51 == io_mem_grant_bits_g_type;
  assign T_2460 = T_2459 ? T_2456 : T_2458;
  assign GEN_52 = {{2'd0}, 2'h0};
  assign T_2461 = GEN_52 == io_mem_grant_bits_g_type;
  assign T_2462 = T_2461 ? 2'h1 : T_2460;
  assign T_2463 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T_2462;
  assign coh_on_grant_state = T_2463;
  assign T_2520 = T_2278 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign coh_on_hit_state = T_2520;
  assign T_2572 = rpq_io_deq_valid == 1'h0;
  assign T_2573 = T_2445 & T_2572;
  assign GEN_1 = T_2573 ? 4'h0 : state;
  assign T_2574 = state == 4'h7;
  assign GEN_2 = T_2574 ? 4'h8 : GEN_1;
  assign T_2575 = state == 4'h6;
  assign T_2576 = T_2575 & io_meta_write_ready;
  assign GEN_3 = T_2576 ? 4'h7 : GEN_2;
  assign T_2577 = state == 4'h5;
  assign T_2578 = T_2577 & refill_done;
  assign GEN_4 = T_2578 ? 4'h6 : GEN_3;
  assign GEN_5 = T_2578 ? coh_on_grant_state : new_coh_state_state;
  assign T_2579 = io_mem_req_ready & io_mem_req_valid;
  assign GEN_6 = T_2579 ? 4'h5 : GEN_4;
  assign T_2580 = state == 4'h3;
  assign T_2581 = T_2580 & io_meta_write_ready;
  assign GEN_7 = T_2581 ? 4'h4 : GEN_6;
  assign T_2582 = state == 4'h2;
  assign T_2583 = T_2582 & io_mem_grant_valid;
  assign GEN_8 = T_2583 ? 4'h3 : GEN_7;
  assign T_2584 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_9 = T_2584 ? 4'h2 : GEN_8;
  assign T_2589 = io_req_sec_val & io_req_sec_rdy;
  assign GEN_10 = cmd_requires_second_acquire ? io_req_bits_cmd : req_cmd;
  assign GEN_11 = T_2589 ? GEN_10 : req_cmd;
  assign T_2607_0 = 2'h2;
  assign T_2607_1 = 2'h3;
  assign T_2609 = T_2607_0 == io_req_bits_old_meta_coh_state;
  assign T_2610 = T_2607_1 == io_req_bits_old_meta_coh_state;
  assign T_2613 = T_2609 | T_2610;
  assign T_2619_0 = 2'h1;
  assign T_2619_1 = 2'h2;
  assign T_2619_2 = 2'h3;
  assign T_2621 = T_2619_0 == io_req_bits_old_meta_coh_state;
  assign T_2622 = T_2619_1 == io_req_bits_old_meta_coh_state;
  assign T_2623 = T_2619_2 == io_req_bits_old_meta_coh_state;
  assign T_2626 = T_2621 | T_2622;
  assign T_2627 = T_2626 | T_2623;
  assign T_2628 = T_2282 ? T_2613 : T_2627;
  assign GEN_12 = T_2628 ? 4'h6 : GEN_9;
  assign GEN_13 = T_2628 ? coh_on_hit_state : GEN_5;
  assign T_2630 = T_2628 == 1'h0;
  assign GEN_14 = T_2630 ? 4'h4 : GEN_12;
  assign GEN_20 = io_req_bits_tag_match ? GEN_14 : GEN_9;
  assign GEN_21 = io_req_bits_tag_match ? GEN_13 : GEN_5;
  assign T_2632 = io_req_bits_tag_match == 1'h0;
  assign T_2638_0 = 2'h3;
  assign T_2640 = T_2638_0 == io_req_bits_old_meta_coh_state;
  assign T_2643 = T_2640 ? 4'h1 : 4'h3;
  assign GEN_23 = T_2632 ? T_2643 : GEN_20;
  assign GEN_24 = T_2436 ? io_req_bits_addr : req_addr;
  assign GEN_25 = T_2436 ? io_req_bits_tag : req_tag;
  assign GEN_26 = T_2436 ? io_req_bits_cmd : GEN_11;
  assign GEN_27 = T_2436 ? io_req_bits_typ : req_typ;
  assign GEN_28 = T_2436 ? io_req_bits_phys : req_phys;
  assign GEN_29 = T_2436 ? io_req_bits_sdq_id : req_sdq_id;
  assign GEN_30 = T_2436 ? io_req_bits_tag_match : req_tag_match;
  assign GEN_31 = T_2436 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign GEN_32 = T_2436 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign GEN_33 = T_2436 ? io_req_bits_way_en : req_way_en;
  assign GEN_39 = T_2436 ? GEN_23 : GEN_9;
  assign GEN_40 = T_2436 ? GEN_21 : GEN_5;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_2682;
  assign fq_io_enq_bits_manager_xact_id = T_2709_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_2709_manager_id;
  assign fq_io_deq_ready = T_2736;
  assign T_2671 = state == 4'h4;
  assign can_finish = T_2447 | T_2671;
  assign GEN_53 = {{1'd0}, 3'h0};
  assign T_2676 = io_mem_grant_bits_g_type == GEN_53;
  assign T_2677 = io_mem_grant_bits_is_builtin_type & T_2676;
  assign T_2679 = T_2677 == 1'h0;
  assign T_2681 = io_mem_grant_valid & T_2679;
  assign T_2682 = T_2681 & refill_done;
  assign T_2709_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign T_2709_manager_id = io_mem_grant_bits_manager_id;
  assign T_2735 = fq_io_deq_valid & can_finish;
  assign T_2736 = io_mem_finish_ready & can_finish;
  assign T_2737 = state != 4'h0;
  assign T_2738 = T_2737 & idx_match;
  assign T_2739 = {req_idx,refill_cnt};
  assign GEN_54 = {{3'd0}, T_2739};
  assign T_2740 = GEN_54 << 3;
  assign T_2741 = req_addr[39:12];
  assign T_2743 = sec_rdy & rpq_io_enq_ready;
  assign GEN_55 = {{1'd0}, 1'h0};
  assign T_2746 = meta_hazard != GEN_55;
  assign GEN_56 = {{1'd0}, 1'h1};
  assign T_2748 = meta_hazard + GEN_56;
  assign T_2749 = T_2748[1:0];
  assign GEN_42 = T_2746 ? T_2749 : meta_hazard;
  assign T_2750 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_43 = T_2750 ? {{1'd0}, 1'h1} : GEN_42;
  assign T_2753 = idx_match == 1'h0;
  assign T_2762 = T_2308 == 1'h0;
  assign T_2764 = meta_hazard == GEN_55;
  assign T_2765 = T_2762 & T_2764;
  assign T_2766 = T_2753 | T_2765;
  assign T_2769 = T_2575 | T_2580;
  assign T_2776_0 = 2'h2;
  assign T_2776_1 = 2'h3;
  assign T_2817_state = 2'h0;
  assign T_2842_state = T_2580 ? T_2817_state : new_coh_state_state;
  assign T_2867 = state == 4'h1;
  assign T_2869 = {req_old_meta_tag,req_idx};
  assign T_2878_0 = 2'h3;
  assign T_2880 = T_2878_0 == req_old_meta_coh_state;
  assign T_2883 = T_2880 ? 3'h0 : 3'h3;
  assign T_2922_addr_beat = {{2'd0}, 1'h0};
  assign T_2922_addr_block = T_2869;
  assign T_2922_client_xact_id = {{1'd0}, 1'h0};
  assign T_2922_voluntary = 1'h1;
  assign T_2922_r_type = T_2883;
  assign T_2922_data = {{63'd0}, 1'h0};
  assign T_2953 = T_2671 & fq_io_enq_ready;
  assign T_2954 = {io_tag,req_idx};
  assign T_2970 = {req_cmd,1'h1};
  assign T_3004_addr_block = T_2954;
  assign T_3004_client_xact_id = {{1'd0}, 1'h0};
  assign T_3004_addr_beat = {{2'd0}, 1'h0};
  assign T_3004_is_builtin_type = 1'h0;
  assign T_3004_a_type = {{2'd0}, T_2293};
  assign T_3004_union = {{6'd0}, T_2970};
  assign T_3004_data = {{63'd0}, 1'h0};
  assign T_3037 = T_2445 & rpq_io_deq_valid;
  assign T_3039 = rpq_io_deq_bits_addr[5:0];
  assign T_3041 = {T_2954,T_3039};
  assign T_3043 = io_meta_read_ready == 1'h0;
  assign GEN_44 = T_3043 ? 1'h0 : T_2448;
  assign GEN_45 = T_3043 ? 5'h5 : rpq_io_deq_bits_cmd;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_16 = {1{$random}};
  state = GEN_16[3:0];
  GEN_17 = {1{$random}};
  new_coh_state_state = GEN_17[1:0];
  GEN_18 = {2{$random}};
  req_addr = GEN_18[39:0];
  GEN_19 = {1{$random}};
  req_tag = GEN_19[8:0];
  GEN_22 = {1{$random}};
  req_cmd = GEN_22[4:0];
  GEN_34 = {1{$random}};
  req_typ = GEN_34[2:0];
  GEN_35 = {1{$random}};
  req_phys = GEN_35[0:0];
  GEN_36 = {1{$random}};
  req_sdq_id = GEN_36[4:0];
  GEN_37 = {1{$random}};
  req_tag_match = GEN_37[0:0];
  GEN_38 = {1{$random}};
  req_old_meta_tag = GEN_38[19:0];
  GEN_41 = {1{$random}};
  req_old_meta_coh_state = GEN_41[1:0];
  GEN_57 = {1{$random}};
  req_way_en = GEN_57[3:0];
  GEN_58 = {1{$random}};
  refill_cnt = GEN_58[2:0];
  GEN_59 = {1{$random}};
  meta_hazard = GEN_59[1:0];
  GEN_60 = {1{$random}};
  GEN_15 = GEN_60[3:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_2436) begin
        if(T_2632) begin
          if(T_2640) begin
            state <= 4'h1;
          end else begin
            state <= 4'h3;
          end
        end else begin
          if(io_req_bits_tag_match) begin
            if(T_2630) begin
              state <= 4'h4;
            end else begin
              if(T_2628) begin
                state <= 4'h6;
              end else begin
                if(T_2584) begin
                  state <= 4'h2;
                end else begin
                  if(T_2583) begin
                    state <= 4'h3;
                  end else begin
                    if(T_2581) begin
                      state <= 4'h4;
                    end else begin
                      if(T_2579) begin
                        state <= 4'h5;
                      end else begin
                        if(T_2578) begin
                          state <= 4'h6;
                        end else begin
                          if(T_2576) begin
                            state <= 4'h7;
                          end else begin
                            if(T_2574) begin
                              state <= 4'h8;
                            end else begin
                              if(T_2573) begin
                                state <= 4'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if(T_2584) begin
              state <= 4'h2;
            end else begin
              if(T_2583) begin
                state <= 4'h3;
              end else begin
                if(T_2581) begin
                  state <= 4'h4;
                end else begin
                  if(T_2579) begin
                    state <= 4'h5;
                  end else begin
                    if(T_2578) begin
                      state <= 4'h6;
                    end else begin
                      if(T_2576) begin
                        state <= 4'h7;
                      end else begin
                        if(T_2574) begin
                          state <= 4'h8;
                        end else begin
                          if(T_2573) begin
                            state <= 4'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if(T_2584) begin
          state <= 4'h2;
        end else begin
          if(T_2583) begin
            state <= 4'h3;
          end else begin
            if(T_2581) begin
              state <= 4'h4;
            end else begin
              if(T_2579) begin
                state <= 4'h5;
              end else begin
                if(T_2578) begin
                  state <= 4'h6;
                end else begin
                  if(T_2576) begin
                    state <= 4'h7;
                  end else begin
                    if(T_2574) begin
                      state <= 4'h8;
                    end else begin
                      if(T_2573) begin
                        state <= 4'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if(reset) begin
      new_coh_state_state <= T_1875_state;
    end else begin
      if(T_2436) begin
        if(io_req_bits_tag_match) begin
          if(T_2628) begin
            new_coh_state_state <= coh_on_hit_state;
          end else begin
            if(T_2578) begin
              new_coh_state_state <= coh_on_grant_state;
            end
          end
        end else begin
          if(T_2578) begin
            new_coh_state_state <= coh_on_grant_state;
          end
        end
      end else begin
        if(T_2578) begin
          new_coh_state_state <= coh_on_grant_state;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_addr <= io_req_bits_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_cmd <= io_req_bits_cmd;
      end else begin
        if(T_2589) begin
          if(cmd_requires_second_acquire) begin
            req_cmd <= io_req_bits_cmd;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_typ <= io_req_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_phys <= io_req_bits_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_sdq_id <= io_req_bits_sdq_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_tag_match <= io_req_bits_tag_match;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_old_meta_tag <= io_req_bits_old_meta_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_way_en <= io_req_bits_way_en;
      end
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      if(T_2350) begin
        refill_cnt <= T_2356;
      end
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else begin
      if(T_2750) begin
        meta_hazard <= {{1'd0}, 1'h1};
      end else begin
        if(T_2746) begin
          meta_hazard <= T_2749;
        end
      end
    end
  end
endmodule
module MSHR_1(
  input   clk,
  input   reset,
  input   io_req_pri_val,
  output  io_req_pri_rdy,
  input   io_req_sec_val,
  output  io_req_sec_rdy,
  input  [39:0] io_req_bits_addr,
  input  [8:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [4:0] io_req_bits_sdq_id,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  output  io_idx_match,
  output [19:0] io_tag,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [11:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [8:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [4:0] io_replay_bits_sdq_id,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy
);
  reg [3:0] state;
  reg [31:0] GEN_16;
  wire [1:0] T_1875_state;
  reg [1:0] new_coh_state_state;
  reg [31:0] GEN_17;
  reg [39:0] req_addr;
  reg [63:0] GEN_18;
  reg [8:0] req_tag;
  reg [31:0] GEN_19;
  reg [4:0] req_cmd;
  reg [31:0] GEN_22;
  reg [2:0] req_typ;
  reg [31:0] GEN_34;
  reg  req_phys;
  reg [31:0] GEN_35;
  reg [4:0] req_sdq_id;
  reg [31:0] GEN_36;
  reg  req_tag_match;
  reg [31:0] GEN_37;
  reg [19:0] req_old_meta_tag;
  reg [31:0] GEN_38;
  reg [1:0] req_old_meta_coh_state;
  reg [31:0] GEN_41;
  reg [3:0] req_way_en;
  reg [31:0] GEN_57;
  wire [5:0] req_idx;
  wire [5:0] T_2271;
  wire  idx_match;
  wire  T_2272;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2278;
  wire  T_2279;
  wire  T_2280;
  wire  T_2281;
  wire  T_2282;
  wire  T_2283;
  wire  T_2284;
  wire  T_2285;
  wire  T_2286;
  wire  T_2287;
  wire  T_2288;
  wire  T_2289;
  wire  T_2290;
  wire  T_2291;
  wire  T_2292;
  wire  T_2293;
  wire  T_2295;
  wire  cmd_requires_second_acquire;
  wire [3:0] states_before_refill_0;
  wire [3:0] states_before_refill_1;
  wire [3:0] states_before_refill_2;
  wire  T_2302;
  wire  T_2303;
  wire  T_2304;
  wire  T_2307;
  wire  T_2308;
  wire [3:0] T_2314_0;
  wire [3:0] T_2314_1;
  wire  T_2316;
  wire  T_2317;
  wire  T_2320;
  wire  T_2322;
  wire  T_2323;
  wire  T_2324;
  wire  sec_rdy;
  wire [2:0] T_2332_0;
  wire [3:0] GEN_46;
  wire  T_2334;
  wire [1:0] T_2342_0;
  wire [1:0] T_2342_1;
  wire [3:0] GEN_47;
  wire  T_2344;
  wire [3:0] GEN_48;
  wire  T_2345;
  wire  T_2348;
  wire  T_2349;
  wire  T_2350;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_58;
  wire  T_2353;
  wire [2:0] GEN_49;
  wire [3:0] T_2355;
  wire [2:0] T_2356;
  wire [2:0] GEN_0;
  wire  refill_count_done;
  wire  T_2358;
  wire  T_2359;
  wire  refill_done;
  wire  rpq_clk;
  wire  rpq_reset;
  wire  rpq_io_enq_ready;
  wire  rpq_io_enq_valid;
  wire [39:0] rpq_io_enq_bits_addr;
  wire [8:0] rpq_io_enq_bits_tag;
  wire [4:0] rpq_io_enq_bits_cmd;
  wire [2:0] rpq_io_enq_bits_typ;
  wire  rpq_io_enq_bits_phys;
  wire [4:0] rpq_io_enq_bits_sdq_id;
  wire  rpq_io_deq_ready;
  wire  rpq_io_deq_valid;
  wire [39:0] rpq_io_deq_bits_addr;
  wire [8:0] rpq_io_deq_bits_tag;
  wire [4:0] rpq_io_deq_bits_cmd;
  wire [2:0] rpq_io_deq_bits_typ;
  wire  rpq_io_deq_bits_phys;
  wire [4:0] rpq_io_deq_bits_sdq_id;
  wire [4:0] rpq_io_count;
  wire  T_2436;
  wire  T_2437;
  wire  T_2438;
  wire  T_2439;
  wire  T_2441;
  wire  T_2443;
  wire  T_2444;
  wire  T_2445;
  wire  T_2446;
  wire  T_2447;
  wire  T_2448;
  wire [1:0] T_2456;
  wire [3:0] GEN_50;
  wire  T_2457;
  wire [1:0] T_2458;
  wire [3:0] GEN_51;
  wire  T_2459;
  wire [1:0] T_2460;
  wire [3:0] GEN_52;
  wire  T_2461;
  wire [1:0] T_2462;
  wire [1:0] T_2463;
  wire [1:0] coh_on_grant_state;
  wire [1:0] T_2520;
  wire [1:0] coh_on_hit_state;
  wire  T_2572;
  wire  T_2573;
  wire [3:0] GEN_1;
  wire  T_2574;
  wire [3:0] GEN_2;
  wire  T_2575;
  wire  T_2576;
  wire [3:0] GEN_3;
  wire  T_2577;
  wire  T_2578;
  wire [3:0] GEN_4;
  wire [1:0] GEN_5;
  wire  T_2579;
  wire [3:0] GEN_6;
  wire  T_2580;
  wire  T_2581;
  wire [3:0] GEN_7;
  wire  T_2582;
  wire  T_2583;
  wire [3:0] GEN_8;
  wire  T_2584;
  wire [3:0] GEN_9;
  wire  T_2589;
  wire [4:0] GEN_10;
  wire [4:0] GEN_11;
  wire [1:0] T_2607_0;
  wire [1:0] T_2607_1;
  wire  T_2609;
  wire  T_2610;
  wire  T_2613;
  wire [1:0] T_2619_0;
  wire [1:0] T_2619_1;
  wire [1:0] T_2619_2;
  wire  T_2621;
  wire  T_2622;
  wire  T_2623;
  wire  T_2626;
  wire  T_2627;
  wire  T_2628;
  wire [3:0] GEN_12;
  wire [1:0] GEN_13;
  wire  T_2630;
  wire [3:0] GEN_14;
  wire [3:0] GEN_20;
  wire [1:0] GEN_21;
  wire  T_2632;
  wire [1:0] T_2638_0;
  wire  T_2640;
  wire [3:0] T_2643;
  wire [3:0] GEN_23;
  wire [39:0] GEN_24;
  wire [8:0] GEN_25;
  wire [4:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [4:0] GEN_29;
  wire  GEN_30;
  wire [19:0] GEN_31;
  wire [1:0] GEN_32;
  wire [3:0] GEN_33;
  wire [3:0] GEN_39;
  wire [1:0] GEN_40;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  wire  T_2671;
  wire  can_finish;
  wire [3:0] GEN_53;
  wire  T_2676;
  wire  T_2677;
  wire  T_2679;
  wire  T_2681;
  wire  T_2682;
  wire [2:0] T_2709_manager_xact_id;
  wire  T_2709_manager_id;
  wire  T_2735;
  wire  T_2736;
  wire  T_2737;
  wire  T_2738;
  wire [8:0] T_2739;
  wire [11:0] GEN_54;
  wire [11:0] T_2740;
  wire [27:0] T_2741;
  wire  T_2743;
  reg [1:0] meta_hazard;
  reg [31:0] GEN_59;
  wire [1:0] GEN_55;
  wire  T_2746;
  wire [1:0] GEN_56;
  wire [2:0] T_2748;
  wire [1:0] T_2749;
  wire [1:0] GEN_42;
  wire  T_2750;
  wire [1:0] GEN_43;
  wire  T_2753;
  wire  T_2762;
  wire  T_2764;
  wire  T_2765;
  wire  T_2766;
  wire  T_2769;
  wire [1:0] T_2776_0;
  wire [1:0] T_2776_1;
  wire [1:0] T_2817_state;
  wire [1:0] T_2842_state;
  wire  T_2867;
  wire [25:0] T_2869;
  wire [1:0] T_2878_0;
  wire  T_2880;
  wire [2:0] T_2883;
  wire [2:0] T_2922_addr_beat;
  wire [25:0] T_2922_addr_block;
  wire [1:0] T_2922_client_xact_id;
  wire  T_2922_voluntary;
  wire [2:0] T_2922_r_type;
  wire [63:0] T_2922_data;
  wire  T_2953;
  wire [25:0] T_2954;
  wire [5:0] T_2970;
  wire [25:0] T_3004_addr_block;
  wire [1:0] T_3004_client_xact_id;
  wire [2:0] T_3004_addr_beat;
  wire  T_3004_is_builtin_type;
  wire [2:0] T_3004_a_type;
  wire [11:0] T_3004_union;
  wire [63:0] T_3004_data;
  wire  T_3037;
  wire [5:0] T_3039;
  wire [31:0] T_3041;
  wire  T_3043;
  wire  GEN_44;
  wire [4:0] GEN_45;
  reg [3:0] GEN_15;
  reg [31:0] GEN_60;
  Queue_1 rpq (
    .clk(rpq_clk),
    .reset(rpq_reset),
    .io_enq_ready(rpq_io_enq_ready),
    .io_enq_valid(rpq_io_enq_valid),
    .io_enq_bits_addr(rpq_io_enq_bits_addr),
    .io_enq_bits_tag(rpq_io_enq_bits_tag),
    .io_enq_bits_cmd(rpq_io_enq_bits_cmd),
    .io_enq_bits_typ(rpq_io_enq_bits_typ),
    .io_enq_bits_phys(rpq_io_enq_bits_phys),
    .io_enq_bits_sdq_id(rpq_io_enq_bits_sdq_id),
    .io_deq_ready(rpq_io_deq_ready),
    .io_deq_valid(rpq_io_deq_valid),
    .io_deq_bits_addr(rpq_io_deq_bits_addr),
    .io_deq_bits_tag(rpq_io_deq_bits_tag),
    .io_deq_bits_cmd(rpq_io_deq_bits_cmd),
    .io_deq_bits_typ(rpq_io_deq_bits_typ),
    .io_deq_bits_phys(rpq_io_deq_bits_phys),
    .io_deq_bits_sdq_id(rpq_io_deq_bits_sdq_id),
    .io_count(rpq_io_count)
  );
  FinishQueue fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_pri_rdy = T_2447;
  assign io_req_sec_rdy = T_2743;
  assign io_idx_match = T_2738;
  assign io_tag = T_2741[19:0];
  assign io_mem_req_valid = T_2953;
  assign io_mem_req_bits_addr_block = T_3004_addr_block;
  assign io_mem_req_bits_client_xact_id = T_3004_client_xact_id;
  assign io_mem_req_bits_addr_beat = T_3004_addr_beat;
  assign io_mem_req_bits_is_builtin_type = T_3004_is_builtin_type;
  assign io_mem_req_bits_a_type = T_3004_a_type;
  assign io_mem_req_bits_union = T_3004_union;
  assign io_mem_req_bits_data = T_3004_data;
  assign io_refill_way_en = req_way_en;
  assign io_refill_addr = T_2740;
  assign io_meta_read_valid = T_2445;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_15;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_write_valid = T_2769;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_data_coh_state = T_2842_state;
  assign io_replay_valid = T_3037;
  assign io_replay_bits_addr = {{8'd0}, T_3041};
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_cmd = GEN_45;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_mem_finish_valid = T_2735;
  assign io_mem_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_wb_req_valid = T_2867;
  assign io_wb_req_bits_addr_beat = T_2922_addr_beat;
  assign io_wb_req_bits_addr_block = T_2922_addr_block;
  assign io_wb_req_bits_client_xact_id = T_2922_client_xact_id;
  assign io_wb_req_bits_voluntary = T_2922_voluntary;
  assign io_wb_req_bits_r_type = T_2922_r_type;
  assign io_wb_req_bits_data = T_2922_data;
  assign io_wb_req_bits_way_en = req_way_en;
  assign io_probe_rdy = T_2766;
  assign T_1875_state = {{1'd0}, 1'h0};
  assign req_idx = req_addr[11:6];
  assign T_2271 = io_req_bits_addr[11:6];
  assign idx_match = req_idx == T_2271;
  assign T_2272 = io_req_bits_cmd == 5'h1;
  assign T_2273 = io_req_bits_cmd == 5'h7;
  assign T_2274 = T_2272 | T_2273;
  assign T_2275 = io_req_bits_cmd[3];
  assign T_2276 = io_req_bits_cmd == 5'h4;
  assign T_2277 = T_2275 | T_2276;
  assign T_2278 = T_2274 | T_2277;
  assign T_2279 = io_req_bits_cmd == 5'h3;
  assign T_2280 = T_2278 | T_2279;
  assign T_2281 = io_req_bits_cmd == 5'h6;
  assign T_2282 = T_2280 | T_2281;
  assign T_2283 = req_cmd == 5'h1;
  assign T_2284 = req_cmd == 5'h7;
  assign T_2285 = T_2283 | T_2284;
  assign T_2286 = req_cmd[3];
  assign T_2287 = req_cmd == 5'h4;
  assign T_2288 = T_2286 | T_2287;
  assign T_2289 = T_2285 | T_2288;
  assign T_2290 = req_cmd == 5'h3;
  assign T_2291 = T_2289 | T_2290;
  assign T_2292 = req_cmd == 5'h6;
  assign T_2293 = T_2291 | T_2292;
  assign T_2295 = T_2293 == 1'h0;
  assign cmd_requires_second_acquire = T_2282 & T_2295;
  assign states_before_refill_0 = 4'h1;
  assign states_before_refill_1 = 4'h2;
  assign states_before_refill_2 = 4'h3;
  assign T_2302 = states_before_refill_0 == state;
  assign T_2303 = states_before_refill_1 == state;
  assign T_2304 = states_before_refill_2 == state;
  assign T_2307 = T_2302 | T_2303;
  assign T_2308 = T_2307 | T_2304;
  assign T_2314_0 = 4'h4;
  assign T_2314_1 = 4'h5;
  assign T_2316 = T_2314_0 == state;
  assign T_2317 = T_2314_1 == state;
  assign T_2320 = T_2316 | T_2317;
  assign T_2322 = cmd_requires_second_acquire == 1'h0;
  assign T_2323 = T_2320 & T_2322;
  assign T_2324 = T_2308 | T_2323;
  assign sec_rdy = idx_match & T_2324;
  assign T_2332_0 = 3'h5;
  assign GEN_46 = {{1'd0}, T_2332_0};
  assign T_2334 = GEN_46 == io_mem_grant_bits_g_type;
  assign T_2342_0 = 2'h0;
  assign T_2342_1 = 2'h1;
  assign GEN_47 = {{2'd0}, T_2342_0};
  assign T_2344 = GEN_47 == io_mem_grant_bits_g_type;
  assign GEN_48 = {{2'd0}, T_2342_1};
  assign T_2345 = GEN_48 == io_mem_grant_bits_g_type;
  assign T_2348 = T_2344 | T_2345;
  assign T_2349 = io_mem_grant_bits_is_builtin_type ? T_2334 : T_2348;
  assign T_2350 = io_mem_grant_valid & T_2349;
  assign T_2353 = refill_cnt == 3'h7;
  assign GEN_49 = {{2'd0}, 1'h1};
  assign T_2355 = refill_cnt + GEN_49;
  assign T_2356 = T_2355[2:0];
  assign GEN_0 = T_2350 ? T_2356 : refill_cnt;
  assign refill_count_done = T_2350 & T_2353;
  assign T_2358 = T_2349 == 1'h0;
  assign T_2359 = T_2358 | refill_count_done;
  assign refill_done = io_mem_grant_valid & T_2359;
  assign rpq_clk = clk;
  assign rpq_reset = reset;
  assign rpq_io_enq_valid = T_2444;
  assign rpq_io_enq_bits_addr = io_req_bits_addr;
  assign rpq_io_enq_bits_tag = io_req_bits_tag;
  assign rpq_io_enq_bits_cmd = io_req_bits_cmd;
  assign rpq_io_enq_bits_typ = io_req_bits_typ;
  assign rpq_io_enq_bits_phys = io_req_bits_phys;
  assign rpq_io_enq_bits_sdq_id = io_req_bits_sdq_id;
  assign rpq_io_deq_ready = GEN_44;
  assign T_2436 = io_req_pri_val & io_req_pri_rdy;
  assign T_2437 = io_req_sec_val & sec_rdy;
  assign T_2438 = T_2436 | T_2437;
  assign T_2439 = io_req_bits_cmd == 5'h2;
  assign T_2441 = T_2439 | T_2279;
  assign T_2443 = T_2441 == 1'h0;
  assign T_2444 = T_2438 & T_2443;
  assign T_2445 = state == 4'h8;
  assign T_2446 = io_replay_ready & T_2445;
  assign T_2447 = state == 4'h0;
  assign T_2448 = T_2446 | T_2447;
  assign T_2456 = T_2289 ? 2'h3 : 2'h2;
  assign GEN_50 = {{2'd0}, 2'h2};
  assign T_2457 = GEN_50 == io_mem_grant_bits_g_type;
  assign T_2458 = T_2457 ? 2'h3 : 2'h0;
  assign GEN_51 = {{2'd0}, 2'h1};
  assign T_2459 = GEN_51 == io_mem_grant_bits_g_type;
  assign T_2460 = T_2459 ? T_2456 : T_2458;
  assign GEN_52 = {{2'd0}, 2'h0};
  assign T_2461 = GEN_52 == io_mem_grant_bits_g_type;
  assign T_2462 = T_2461 ? 2'h1 : T_2460;
  assign T_2463 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T_2462;
  assign coh_on_grant_state = T_2463;
  assign T_2520 = T_2278 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign coh_on_hit_state = T_2520;
  assign T_2572 = rpq_io_deq_valid == 1'h0;
  assign T_2573 = T_2445 & T_2572;
  assign GEN_1 = T_2573 ? 4'h0 : state;
  assign T_2574 = state == 4'h7;
  assign GEN_2 = T_2574 ? 4'h8 : GEN_1;
  assign T_2575 = state == 4'h6;
  assign T_2576 = T_2575 & io_meta_write_ready;
  assign GEN_3 = T_2576 ? 4'h7 : GEN_2;
  assign T_2577 = state == 4'h5;
  assign T_2578 = T_2577 & refill_done;
  assign GEN_4 = T_2578 ? 4'h6 : GEN_3;
  assign GEN_5 = T_2578 ? coh_on_grant_state : new_coh_state_state;
  assign T_2579 = io_mem_req_ready & io_mem_req_valid;
  assign GEN_6 = T_2579 ? 4'h5 : GEN_4;
  assign T_2580 = state == 4'h3;
  assign T_2581 = T_2580 & io_meta_write_ready;
  assign GEN_7 = T_2581 ? 4'h4 : GEN_6;
  assign T_2582 = state == 4'h2;
  assign T_2583 = T_2582 & io_mem_grant_valid;
  assign GEN_8 = T_2583 ? 4'h3 : GEN_7;
  assign T_2584 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_9 = T_2584 ? 4'h2 : GEN_8;
  assign T_2589 = io_req_sec_val & io_req_sec_rdy;
  assign GEN_10 = cmd_requires_second_acquire ? io_req_bits_cmd : req_cmd;
  assign GEN_11 = T_2589 ? GEN_10 : req_cmd;
  assign T_2607_0 = 2'h2;
  assign T_2607_1 = 2'h3;
  assign T_2609 = T_2607_0 == io_req_bits_old_meta_coh_state;
  assign T_2610 = T_2607_1 == io_req_bits_old_meta_coh_state;
  assign T_2613 = T_2609 | T_2610;
  assign T_2619_0 = 2'h1;
  assign T_2619_1 = 2'h2;
  assign T_2619_2 = 2'h3;
  assign T_2621 = T_2619_0 == io_req_bits_old_meta_coh_state;
  assign T_2622 = T_2619_1 == io_req_bits_old_meta_coh_state;
  assign T_2623 = T_2619_2 == io_req_bits_old_meta_coh_state;
  assign T_2626 = T_2621 | T_2622;
  assign T_2627 = T_2626 | T_2623;
  assign T_2628 = T_2282 ? T_2613 : T_2627;
  assign GEN_12 = T_2628 ? 4'h6 : GEN_9;
  assign GEN_13 = T_2628 ? coh_on_hit_state : GEN_5;
  assign T_2630 = T_2628 == 1'h0;
  assign GEN_14 = T_2630 ? 4'h4 : GEN_12;
  assign GEN_20 = io_req_bits_tag_match ? GEN_14 : GEN_9;
  assign GEN_21 = io_req_bits_tag_match ? GEN_13 : GEN_5;
  assign T_2632 = io_req_bits_tag_match == 1'h0;
  assign T_2638_0 = 2'h3;
  assign T_2640 = T_2638_0 == io_req_bits_old_meta_coh_state;
  assign T_2643 = T_2640 ? 4'h1 : 4'h3;
  assign GEN_23 = T_2632 ? T_2643 : GEN_20;
  assign GEN_24 = T_2436 ? io_req_bits_addr : req_addr;
  assign GEN_25 = T_2436 ? io_req_bits_tag : req_tag;
  assign GEN_26 = T_2436 ? io_req_bits_cmd : GEN_11;
  assign GEN_27 = T_2436 ? io_req_bits_typ : req_typ;
  assign GEN_28 = T_2436 ? io_req_bits_phys : req_phys;
  assign GEN_29 = T_2436 ? io_req_bits_sdq_id : req_sdq_id;
  assign GEN_30 = T_2436 ? io_req_bits_tag_match : req_tag_match;
  assign GEN_31 = T_2436 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign GEN_32 = T_2436 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign GEN_33 = T_2436 ? io_req_bits_way_en : req_way_en;
  assign GEN_39 = T_2436 ? GEN_23 : GEN_9;
  assign GEN_40 = T_2436 ? GEN_21 : GEN_5;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_2682;
  assign fq_io_enq_bits_manager_xact_id = T_2709_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_2709_manager_id;
  assign fq_io_deq_ready = T_2736;
  assign T_2671 = state == 4'h4;
  assign can_finish = T_2447 | T_2671;
  assign GEN_53 = {{1'd0}, 3'h0};
  assign T_2676 = io_mem_grant_bits_g_type == GEN_53;
  assign T_2677 = io_mem_grant_bits_is_builtin_type & T_2676;
  assign T_2679 = T_2677 == 1'h0;
  assign T_2681 = io_mem_grant_valid & T_2679;
  assign T_2682 = T_2681 & refill_done;
  assign T_2709_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign T_2709_manager_id = io_mem_grant_bits_manager_id;
  assign T_2735 = fq_io_deq_valid & can_finish;
  assign T_2736 = io_mem_finish_ready & can_finish;
  assign T_2737 = state != 4'h0;
  assign T_2738 = T_2737 & idx_match;
  assign T_2739 = {req_idx,refill_cnt};
  assign GEN_54 = {{3'd0}, T_2739};
  assign T_2740 = GEN_54 << 3;
  assign T_2741 = req_addr[39:12];
  assign T_2743 = sec_rdy & rpq_io_enq_ready;
  assign GEN_55 = {{1'd0}, 1'h0};
  assign T_2746 = meta_hazard != GEN_55;
  assign GEN_56 = {{1'd0}, 1'h1};
  assign T_2748 = meta_hazard + GEN_56;
  assign T_2749 = T_2748[1:0];
  assign GEN_42 = T_2746 ? T_2749 : meta_hazard;
  assign T_2750 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_43 = T_2750 ? {{1'd0}, 1'h1} : GEN_42;
  assign T_2753 = idx_match == 1'h0;
  assign T_2762 = T_2308 == 1'h0;
  assign T_2764 = meta_hazard == GEN_55;
  assign T_2765 = T_2762 & T_2764;
  assign T_2766 = T_2753 | T_2765;
  assign T_2769 = T_2575 | T_2580;
  assign T_2776_0 = 2'h2;
  assign T_2776_1 = 2'h3;
  assign T_2817_state = 2'h0;
  assign T_2842_state = T_2580 ? T_2817_state : new_coh_state_state;
  assign T_2867 = state == 4'h1;
  assign T_2869 = {req_old_meta_tag,req_idx};
  assign T_2878_0 = 2'h3;
  assign T_2880 = T_2878_0 == req_old_meta_coh_state;
  assign T_2883 = T_2880 ? 3'h0 : 3'h3;
  assign T_2922_addr_beat = {{2'd0}, 1'h0};
  assign T_2922_addr_block = T_2869;
  assign T_2922_client_xact_id = {{1'd0}, 1'h1};
  assign T_2922_voluntary = 1'h1;
  assign T_2922_r_type = T_2883;
  assign T_2922_data = {{63'd0}, 1'h0};
  assign T_2953 = T_2671 & fq_io_enq_ready;
  assign T_2954 = {io_tag,req_idx};
  assign T_2970 = {req_cmd,1'h1};
  assign T_3004_addr_block = T_2954;
  assign T_3004_client_xact_id = {{1'd0}, 1'h1};
  assign T_3004_addr_beat = {{2'd0}, 1'h0};
  assign T_3004_is_builtin_type = 1'h0;
  assign T_3004_a_type = {{2'd0}, T_2293};
  assign T_3004_union = {{6'd0}, T_2970};
  assign T_3004_data = {{63'd0}, 1'h0};
  assign T_3037 = T_2445 & rpq_io_deq_valid;
  assign T_3039 = rpq_io_deq_bits_addr[5:0];
  assign T_3041 = {T_2954,T_3039};
  assign T_3043 = io_meta_read_ready == 1'h0;
  assign GEN_44 = T_3043 ? 1'h0 : T_2448;
  assign GEN_45 = T_3043 ? 5'h5 : rpq_io_deq_bits_cmd;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_16 = {1{$random}};
  state = GEN_16[3:0];
  GEN_17 = {1{$random}};
  new_coh_state_state = GEN_17[1:0];
  GEN_18 = {2{$random}};
  req_addr = GEN_18[39:0];
  GEN_19 = {1{$random}};
  req_tag = GEN_19[8:0];
  GEN_22 = {1{$random}};
  req_cmd = GEN_22[4:0];
  GEN_34 = {1{$random}};
  req_typ = GEN_34[2:0];
  GEN_35 = {1{$random}};
  req_phys = GEN_35[0:0];
  GEN_36 = {1{$random}};
  req_sdq_id = GEN_36[4:0];
  GEN_37 = {1{$random}};
  req_tag_match = GEN_37[0:0];
  GEN_38 = {1{$random}};
  req_old_meta_tag = GEN_38[19:0];
  GEN_41 = {1{$random}};
  req_old_meta_coh_state = GEN_41[1:0];
  GEN_57 = {1{$random}};
  req_way_en = GEN_57[3:0];
  GEN_58 = {1{$random}};
  refill_cnt = GEN_58[2:0];
  GEN_59 = {1{$random}};
  meta_hazard = GEN_59[1:0];
  GEN_60 = {1{$random}};
  GEN_15 = GEN_60[3:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_2436) begin
        if(T_2632) begin
          if(T_2640) begin
            state <= 4'h1;
          end else begin
            state <= 4'h3;
          end
        end else begin
          if(io_req_bits_tag_match) begin
            if(T_2630) begin
              state <= 4'h4;
            end else begin
              if(T_2628) begin
                state <= 4'h6;
              end else begin
                if(T_2584) begin
                  state <= 4'h2;
                end else begin
                  if(T_2583) begin
                    state <= 4'h3;
                  end else begin
                    if(T_2581) begin
                      state <= 4'h4;
                    end else begin
                      if(T_2579) begin
                        state <= 4'h5;
                      end else begin
                        if(T_2578) begin
                          state <= 4'h6;
                        end else begin
                          if(T_2576) begin
                            state <= 4'h7;
                          end else begin
                            if(T_2574) begin
                              state <= 4'h8;
                            end else begin
                              if(T_2573) begin
                                state <= 4'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if(T_2584) begin
              state <= 4'h2;
            end else begin
              if(T_2583) begin
                state <= 4'h3;
              end else begin
                if(T_2581) begin
                  state <= 4'h4;
                end else begin
                  if(T_2579) begin
                    state <= 4'h5;
                  end else begin
                    if(T_2578) begin
                      state <= 4'h6;
                    end else begin
                      if(T_2576) begin
                        state <= 4'h7;
                      end else begin
                        if(T_2574) begin
                          state <= 4'h8;
                        end else begin
                          if(T_2573) begin
                            state <= 4'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if(T_2584) begin
          state <= 4'h2;
        end else begin
          if(T_2583) begin
            state <= 4'h3;
          end else begin
            if(T_2581) begin
              state <= 4'h4;
            end else begin
              if(T_2579) begin
                state <= 4'h5;
              end else begin
                if(T_2578) begin
                  state <= 4'h6;
                end else begin
                  if(T_2576) begin
                    state <= 4'h7;
                  end else begin
                    if(T_2574) begin
                      state <= 4'h8;
                    end else begin
                      if(T_2573) begin
                        state <= 4'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if(reset) begin
      new_coh_state_state <= T_1875_state;
    end else begin
      if(T_2436) begin
        if(io_req_bits_tag_match) begin
          if(T_2628) begin
            new_coh_state_state <= coh_on_hit_state;
          end else begin
            if(T_2578) begin
              new_coh_state_state <= coh_on_grant_state;
            end
          end
        end else begin
          if(T_2578) begin
            new_coh_state_state <= coh_on_grant_state;
          end
        end
      end else begin
        if(T_2578) begin
          new_coh_state_state <= coh_on_grant_state;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_addr <= io_req_bits_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_cmd <= io_req_bits_cmd;
      end else begin
        if(T_2589) begin
          if(cmd_requires_second_acquire) begin
            req_cmd <= io_req_bits_cmd;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_typ <= io_req_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_phys <= io_req_bits_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_sdq_id <= io_req_bits_sdq_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_tag_match <= io_req_bits_tag_match;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_old_meta_tag <= io_req_bits_old_meta_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2436) begin
        req_way_en <= io_req_bits_way_en;
      end
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      if(T_2350) begin
        refill_cnt <= T_2356;
      end
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else begin
      if(T_2750) begin
        meta_hazard <= {{1'd0}, 1'h1};
      end else begin
        if(T_2746) begin
          meta_hazard <= T_2749;
        end
      end
    end
  end
endmodule
module Arbiter_6(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits,
  input   io_out_ready,
  output  io_out_valid,
  output  io_out_bits,
  output  io_chosen
);
  assign io_in_0_ready = io_out_ready;
  assign io_out_valid = io_in_0_valid;
  assign io_out_bits = io_in_0_bits;
  assign io_chosen = 1'h0;
endmodule
module Arbiter_7(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [8:0] io_in_0_bits_tag,
  input  [4:0] io_in_0_bits_cmd,
  input  [2:0] io_in_0_bits_typ,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_replay,
  input   io_in_0_bits_has_data,
  input  [63:0] io_in_0_bits_data_word_bypass,
  input  [63:0] io_in_0_bits_store_data,
  input   io_out_ready,
  output  io_out_valid,
  output [39:0] io_out_bits_addr,
  output [8:0] io_out_bits_tag,
  output [4:0] io_out_bits_cmd,
  output [2:0] io_out_bits_typ,
  output [63:0] io_out_bits_data,
  output  io_out_bits_replay,
  output  io_out_bits_has_data,
  output [63:0] io_out_bits_data_word_bypass,
  output [63:0] io_out_bits_store_data,
  output  io_chosen
);
  assign io_in_0_ready = io_out_ready;
  assign io_out_valid = io_in_0_valid;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_bits_cmd = io_in_0_bits_cmd;
  assign io_out_bits_typ = io_in_0_bits_typ;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_bits_replay = io_in_0_bits_replay;
  assign io_out_bits_has_data = io_in_0_bits_has_data;
  assign io_out_bits_data_word_bypass = io_in_0_bits_data_word_bypass;
  assign io_out_bits_store_data = io_in_0_bits_store_data;
  assign io_chosen = 1'h0;
endmodule
module IOMSHR(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [39:0] io_req_bits_addr,
  input  [8:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [63:0] io_req_bits_data,
  input   io_acquire_ready,
  output  io_acquire_valid,
  output [25:0] io_acquire_bits_addr_block,
  output [1:0] io_acquire_bits_client_xact_id,
  output [2:0] io_acquire_bits_addr_beat,
  output  io_acquire_bits_is_builtin_type,
  output [2:0] io_acquire_bits_a_type,
  output [11:0] io_acquire_bits_union,
  output [63:0] io_acquire_bits_data,
  input   io_grant_valid,
  input  [2:0] io_grant_bits_addr_beat,
  input  [1:0] io_grant_bits_client_xact_id,
  input  [2:0] io_grant_bits_manager_xact_id,
  input   io_grant_bits_is_builtin_type,
  input  [3:0] io_grant_bits_g_type,
  input  [63:0] io_grant_bits_data,
  input   io_grant_bits_manager_id,
  input   io_finish_ready,
  output  io_finish_valid,
  output [2:0] io_finish_bits_manager_xact_id,
  output  io_finish_bits_manager_id,
  input   io_resp_ready,
  output  io_resp_valid,
  output [39:0] io_resp_bits_addr,
  output [8:0] io_resp_bits_tag,
  output [4:0] io_resp_bits_cmd,
  output [2:0] io_resp_bits_typ,
  output [63:0] io_resp_bits_data,
  output  io_resp_bits_replay,
  output  io_resp_bits_has_data,
  output [63:0] io_resp_bits_data_word_bypass,
  output [63:0] io_resp_bits_store_data,
  output  io_replay_next
);
  reg [39:0] req_addr;
  reg [63:0] GEN_22;
  reg [8:0] req_tag;
  reg [31:0] GEN_24;
  reg [4:0] req_cmd;
  reg [31:0] GEN_27;
  reg [2:0] req_typ;
  reg [31:0] GEN_28;
  reg  req_phys;
  reg [31:0] GEN_29;
  reg [63:0] req_data;
  reg [63:0] GEN_30;
  wire  req_cmd_sc;
  reg [63:0] grant_word;
  reg [63:0] GEN_31;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  reg [2:0] state;
  reg [31:0] GEN_32;
  wire  T_1211;
  wire [3:0] GEN_13;
  wire  T_1216;
  wire  T_1217;
  wire  T_1219;
  wire  T_1221;
  wire [2:0] T_1248_manager_xact_id;
  wire  T_1248_manager_id;
  wire  T_1274;
  wire  T_1275;
  wire  T_1277;
  wire [1:0] T_1278;
  wire [2:0] T_1280;
  wire  GEN_14;
  wire [2:0] GEN_15;
  wire  T_1282;
  wire  T_1284;
  wire [1:0] GEN_16;
  wire  T_1288;
  wire  T_1292;
  wire  T_1295;
  wire [1:0] T_1296;
  wire  T_1297;
  wire [1:0] T_1299;
  wire  T_1301;
  wire [1:0] T_1304;
  wire [1:0] T_1305;
  wire [1:0] T_1308;
  wire [3:0] T_1309;
  wire  T_1310;
  wire [3:0] T_1312;
  wire  T_1314;
  wire [3:0] T_1317;
  wire [3:0] T_1318;
  wire [3:0] T_1321;
  wire [7:0] T_1322;
  wire [22:0] GEN_17;
  wire [22:0] beat_mask;
  wire [1:0] GEN_18;
  wire  T_1327;
  wire [7:0] T_1328;
  wire [15:0] T_1329;
  wire [31:0] T_1330;
  wire [63:0] T_1331;
  wire  T_1333;
  wire [15:0] T_1334;
  wire [31:0] T_1335;
  wire [63:0] T_1336;
  wire  T_1338;
  wire [31:0] T_1339;
  wire [63:0] T_1340;
  wire [63:0] T_1341;
  wire [63:0] T_1342;
  wire [63:0] beat_data;
  wire [25:0] addr_block;
  wire [2:0] addr_beat;
  wire [2:0] addr_byte;
  wire [5:0] T_1387;
  wire [11:0] T_1388;
  wire [25:0] get_acquire_addr_block;
  wire [1:0] get_acquire_client_xact_id;
  wire [2:0] get_acquire_addr_beat;
  wire  get_acquire_is_builtin_type;
  wire [2:0] get_acquire_a_type;
  wire [11:0] get_acquire_union;
  wire [63:0] get_acquire_data;
  wire [22:0] GEN_20;
  wire [22:0] T_1518;
  wire [7:0] T_1519;
  wire [8:0] T_1529;
  wire [11:0] T_1549;
  wire [25:0] put_acquire_addr_block;
  wire [1:0] put_acquire_client_xact_id;
  wire [2:0] put_acquire_addr_beat;
  wire  put_acquire_is_builtin_type;
  wire [2:0] put_acquire_a_type;
  wire [11:0] put_acquire_union;
  wire [63:0] put_acquire_data;
  wire [5:0] T_1657;
  wire [11:0] T_1659;
  wire [25:0] putAtomic_acquire_addr_block;
  wire [1:0] putAtomic_acquire_client_xact_id;
  wire [2:0] putAtomic_acquire_addr_beat;
  wire  putAtomic_acquire_is_builtin_type;
  wire [2:0] putAtomic_acquire_a_type;
  wire [11:0] putAtomic_acquire_union;
  wire [63:0] putAtomic_acquire_data;
  wire  T_1750;
  wire  T_1751;
  wire  T_1752;
  wire  T_1753;
  wire  T_1754;
  wire  T_1755;
  wire  T_1756;
  wire  T_1758;
  wire  T_1762;
  wire [25:0] T_1763_addr_block;
  wire [1:0] T_1763_client_xact_id;
  wire [2:0] T_1763_addr_beat;
  wire  T_1763_is_builtin_type;
  wire [2:0] T_1763_a_type;
  wire [11:0] T_1763_union;
  wire [63:0] T_1763_data;
  wire [25:0] T_1794_addr_block;
  wire [1:0] T_1794_client_xact_id;
  wire [2:0] T_1794_addr_beat;
  wire  T_1794_is_builtin_type;
  wire [2:0] T_1794_a_type;
  wire [11:0] T_1794_union;
  wire [63:0] T_1794_data;
  wire  T_1825;
  wire  T_1827;
  wire  T_1828;
  wire  T_1829;
  wire  T_1830;
  wire [31:0] T_1841;
  wire [31:0] T_1842;
  wire [31:0] T_1843;
  wire  T_1851;
  wire  T_1852;
  wire [31:0] GEN_21;
  wire [32:0] T_1854;
  wire [31:0] T_1855;
  wire [31:0] T_1857;
  wire [63:0] T_1858;
  wire [15:0] T_1860;
  wire [15:0] T_1861;
  wire [15:0] T_1862;
  wire  T_1870;
  wire  T_1871;
  wire [47:0] GEN_23;
  wire [48:0] T_1873;
  wire [47:0] T_1874;
  wire [47:0] T_1875;
  wire [47:0] T_1876;
  wire [63:0] T_1877;
  wire [7:0] T_1879;
  wire [7:0] T_1880;
  wire [7:0] T_1881;
  wire [7:0] T_1885;
  wire  T_1888;
  wire  T_1889;
  wire  T_1890;
  wire [55:0] GEN_25;
  wire [56:0] T_1892;
  wire [55:0] T_1893;
  wire [55:0] T_1894;
  wire [55:0] T_1895;
  wire [63:0] T_1896;
  wire [63:0] GEN_26;
  wire [63:0] T_1897;
  wire  T_1899;
  wire [39:0] GEN_0;
  wire [8:0] GEN_1;
  wire [4:0] GEN_2;
  wire [2:0] GEN_3;
  wire  GEN_4;
  wire [63:0] GEN_5;
  wire [2:0] GEN_6;
  wire  T_1900;
  wire [2:0] GEN_7;
  wire  T_1902;
  wire [63:0] T_1915;
  wire [63:0] GEN_8;
  wire [2:0] GEN_9;
  wire [63:0] GEN_10;
  wire  T_1917;
  wire [2:0] GEN_11;
  wire  T_1918;
  wire [2:0] GEN_12;
  reg [63:0] GEN_19;
  reg [63:0] GEN_33;
  FinishQueue fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_ready = T_1211;
  assign io_acquire_valid = T_1750;
  assign io_acquire_bits_addr_block = T_1794_addr_block;
  assign io_acquire_bits_client_xact_id = T_1794_client_xact_id;
  assign io_acquire_bits_addr_beat = T_1794_addr_beat;
  assign io_acquire_bits_is_builtin_type = T_1794_is_builtin_type;
  assign io_acquire_bits_a_type = T_1794_a_type;
  assign io_acquire_bits_union = T_1794_union;
  assign io_acquire_bits_data = T_1794_data;
  assign io_finish_valid = T_1275;
  assign io_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_resp_valid = T_1830;
  assign io_resp_bits_addr = req_addr;
  assign io_resp_bits_tag = req_tag;
  assign io_resp_bits_cmd = req_cmd;
  assign io_resp_bits_typ = req_typ;
  assign io_resp_bits_data = T_1897;
  assign io_resp_bits_replay = 1'h1;
  assign io_resp_bits_has_data = T_1762;
  assign io_resp_bits_data_word_bypass = GEN_19;
  assign io_resp_bits_store_data = req_data;
  assign io_replay_next = T_1829;
  assign req_cmd_sc = req_cmd == 5'h7;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_1221;
  assign fq_io_enq_bits_manager_xact_id = T_1248_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_1248_manager_id;
  assign fq_io_deq_ready = T_1277;
  assign T_1211 = state == 3'h0;
  assign GEN_13 = {{1'd0}, 3'h0};
  assign T_1216 = io_grant_bits_g_type == GEN_13;
  assign T_1217 = io_grant_bits_is_builtin_type & T_1216;
  assign T_1219 = T_1217 == 1'h0;
  assign T_1221 = io_grant_valid & T_1219;
  assign T_1248_manager_xact_id = io_grant_bits_manager_xact_id;
  assign T_1248_manager_id = io_grant_bits_manager_id;
  assign T_1274 = state == 3'h4;
  assign T_1275 = fq_io_deq_valid & T_1274;
  assign T_1277 = io_finish_ready & T_1274;
  assign T_1278 = req_typ[1:0];
  assign T_1280 = $signed(req_typ);
  assign GEN_14 = $signed(1'h0);
  assign GEN_15 = {3{GEN_14}};
  assign T_1282 = $signed(T_1280) >= $signed(GEN_15);
  assign T_1284 = req_addr[0];
  assign GEN_16 = {{1'd0}, 1'h1};
  assign T_1288 = T_1278 >= GEN_16;
  assign T_1292 = T_1284 | T_1288;
  assign T_1295 = T_1284 ? 1'h0 : 1'h1;
  assign T_1296 = {T_1292,T_1295};
  assign T_1297 = req_addr[1];
  assign T_1299 = T_1297 ? T_1296 : {{1'd0}, 1'h0};
  assign T_1301 = T_1278 >= 2'h2;
  assign T_1304 = T_1301 ? 2'h3 : {{1'd0}, 1'h0};
  assign T_1305 = T_1299 | T_1304;
  assign T_1308 = T_1297 ? {{1'd0}, 1'h0} : T_1296;
  assign T_1309 = {T_1305,T_1308};
  assign T_1310 = req_addr[2];
  assign T_1312 = T_1310 ? T_1309 : {{3'd0}, 1'h0};
  assign T_1314 = T_1278 >= 2'h3;
  assign T_1317 = T_1314 ? 4'hf : {{3'd0}, 1'h0};
  assign T_1318 = T_1312 | T_1317;
  assign T_1321 = T_1310 ? {{3'd0}, 1'h0} : T_1309;
  assign T_1322 = {T_1318,T_1321};
  assign GEN_17 = {{15'd0}, T_1322};
  assign beat_mask = GEN_17 << 4'h0;
  assign GEN_18 = {{1'd0}, 1'h0};
  assign T_1327 = T_1278 == GEN_18;
  assign T_1328 = req_data[7:0];
  assign T_1329 = {T_1328,T_1328};
  assign T_1330 = {T_1329,T_1329};
  assign T_1331 = {T_1330,T_1330};
  assign T_1333 = T_1278 == GEN_16;
  assign T_1334 = req_data[15:0];
  assign T_1335 = {T_1334,T_1334};
  assign T_1336 = {T_1335,T_1335};
  assign T_1338 = T_1278 == 2'h2;
  assign T_1339 = req_data[31:0];
  assign T_1340 = {T_1339,T_1339};
  assign T_1341 = T_1338 ? T_1340 : req_data;
  assign T_1342 = T_1333 ? T_1336 : T_1341;
  assign beat_data = T_1327 ? T_1331 : T_1342;
  assign addr_block = req_addr[31:6];
  assign addr_beat = req_addr[5:3];
  assign addr_byte = req_addr[2:0];
  assign T_1387 = {addr_byte,req_typ};
  assign T_1388 = {T_1387,6'h0};
  assign get_acquire_addr_block = addr_block;
  assign get_acquire_client_xact_id = 2'h2;
  assign get_acquire_addr_beat = addr_beat;
  assign get_acquire_is_builtin_type = 1'h1;
  assign get_acquire_a_type = 3'h0;
  assign get_acquire_union = T_1388;
  assign get_acquire_data = {{63'd0}, 1'h0};
  assign GEN_20 = {{15'd0}, 8'h0};
  assign T_1518 = GEN_20 | beat_mask;
  assign T_1519 = T_1518[7:0];
  assign T_1529 = {T_1519,1'h0};
  assign T_1549 = 1'h1 ? {{3'd0}, T_1529} : 12'h0;
  assign put_acquire_addr_block = addr_block;
  assign put_acquire_client_xact_id = 2'h2;
  assign put_acquire_addr_beat = addr_beat;
  assign put_acquire_is_builtin_type = 1'h1;
  assign put_acquire_a_type = 3'h2;
  assign put_acquire_union = T_1549;
  assign put_acquire_data = beat_data;
  assign T_1657 = {req_cmd,1'h1};
  assign T_1659 = {T_1387,T_1657};
  assign putAtomic_acquire_addr_block = addr_block;
  assign putAtomic_acquire_client_xact_id = 2'h2;
  assign putAtomic_acquire_addr_beat = addr_beat;
  assign putAtomic_acquire_is_builtin_type = 1'h1;
  assign putAtomic_acquire_a_type = 3'h4;
  assign putAtomic_acquire_union = T_1659;
  assign putAtomic_acquire_data = beat_data;
  assign T_1750 = state == 3'h1;
  assign T_1751 = req_cmd[3];
  assign T_1752 = req_cmd == 5'h4;
  assign T_1753 = T_1751 | T_1752;
  assign T_1754 = req_cmd == 5'h0;
  assign T_1755 = req_cmd == 5'h6;
  assign T_1756 = T_1754 | T_1755;
  assign T_1758 = T_1756 | req_cmd_sc;
  assign T_1762 = T_1758 | T_1753;
  assign T_1763_addr_block = T_1762 ? get_acquire_addr_block : put_acquire_addr_block;
  assign T_1763_client_xact_id = T_1762 ? get_acquire_client_xact_id : put_acquire_client_xact_id;
  assign T_1763_addr_beat = T_1762 ? get_acquire_addr_beat : put_acquire_addr_beat;
  assign T_1763_is_builtin_type = T_1762 ? get_acquire_is_builtin_type : put_acquire_is_builtin_type;
  assign T_1763_a_type = T_1762 ? get_acquire_a_type : put_acquire_a_type;
  assign T_1763_union = T_1762 ? get_acquire_union : put_acquire_union;
  assign T_1763_data = T_1762 ? get_acquire_data : put_acquire_data;
  assign T_1794_addr_block = T_1753 ? putAtomic_acquire_addr_block : T_1763_addr_block;
  assign T_1794_client_xact_id = T_1753 ? putAtomic_acquire_client_xact_id : T_1763_client_xact_id;
  assign T_1794_addr_beat = T_1753 ? putAtomic_acquire_addr_beat : T_1763_addr_beat;
  assign T_1794_is_builtin_type = T_1753 ? putAtomic_acquire_is_builtin_type : T_1763_is_builtin_type;
  assign T_1794_a_type = T_1753 ? putAtomic_acquire_a_type : T_1763_a_type;
  assign T_1794_union = T_1753 ? putAtomic_acquire_union : T_1763_union;
  assign T_1794_data = T_1753 ? putAtomic_acquire_data : T_1763_data;
  assign T_1825 = state == 3'h2;
  assign T_1827 = io_resp_ready == 1'h0;
  assign T_1828 = io_resp_valid & T_1827;
  assign T_1829 = T_1825 | T_1828;
  assign T_1830 = state == 3'h3;
  assign T_1841 = grant_word[63:32];
  assign T_1842 = grant_word[31:0];
  assign T_1843 = T_1310 ? T_1841 : T_1842;
  assign T_1851 = T_1843[31];
  assign T_1852 = T_1282 & T_1851;
  assign GEN_21 = {{31'd0}, T_1852};
  assign T_1854 = 32'h0 - GEN_21;
  assign T_1855 = T_1854[31:0];
  assign T_1857 = T_1338 ? T_1855 : T_1841;
  assign T_1858 = {T_1857,T_1843};
  assign T_1860 = T_1858[31:16];
  assign T_1861 = T_1858[15:0];
  assign T_1862 = T_1297 ? T_1860 : T_1861;
  assign T_1870 = T_1862[15];
  assign T_1871 = T_1282 & T_1870;
  assign GEN_23 = {{47'd0}, T_1871};
  assign T_1873 = 48'h0 - GEN_23;
  assign T_1874 = T_1873[47:0];
  assign T_1875 = T_1858[63:16];
  assign T_1876 = T_1333 ? T_1874 : T_1875;
  assign T_1877 = {T_1876,T_1862};
  assign T_1879 = T_1877[15:8];
  assign T_1880 = T_1877[7:0];
  assign T_1881 = T_1284 ? T_1879 : T_1880;
  assign T_1885 = req_cmd_sc ? {{7'd0}, 1'h0} : T_1881;
  assign T_1888 = T_1327 | req_cmd_sc;
  assign T_1889 = T_1885[7];
  assign T_1890 = T_1282 & T_1889;
  assign GEN_25 = {{55'd0}, T_1890};
  assign T_1892 = 56'h0 - GEN_25;
  assign T_1893 = T_1892[55:0];
  assign T_1894 = T_1877[63:8];
  assign T_1895 = T_1888 ? T_1893 : T_1894;
  assign T_1896 = {T_1895,T_1885};
  assign GEN_26 = {{63'd0}, req_cmd_sc};
  assign T_1897 = T_1896 | GEN_26;
  assign T_1899 = io_req_ready & io_req_valid;
  assign GEN_0 = T_1899 ? io_req_bits_addr : req_addr;
  assign GEN_1 = T_1899 ? io_req_bits_tag : req_tag;
  assign GEN_2 = T_1899 ? io_req_bits_cmd : req_cmd;
  assign GEN_3 = T_1899 ? io_req_bits_typ : req_typ;
  assign GEN_4 = T_1899 ? io_req_bits_phys : req_phys;
  assign GEN_5 = T_1899 ? io_req_bits_data : req_data;
  assign GEN_6 = T_1899 ? 3'h1 : state;
  assign T_1900 = io_acquire_ready & io_acquire_valid;
  assign GEN_7 = T_1900 ? 3'h2 : GEN_6;
  assign T_1902 = T_1825 & io_grant_valid;
  assign T_1915 = io_grant_bits_data >> 7'h0;
  assign GEN_8 = T_1762 ? T_1915 : grant_word;
  assign GEN_9 = T_1902 ? 3'h3 : GEN_7;
  assign GEN_10 = T_1902 ? GEN_8 : grant_word;
  assign T_1917 = io_resp_ready & io_resp_valid;
  assign GEN_11 = T_1917 ? 3'h4 : GEN_9;
  assign T_1918 = io_finish_ready & io_finish_valid;
  assign GEN_12 = T_1918 ? 3'h0 : GEN_11;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_22 = {2{$random}};
  req_addr = GEN_22[39:0];
  GEN_24 = {1{$random}};
  req_tag = GEN_24[8:0];
  GEN_27 = {1{$random}};
  req_cmd = GEN_27[4:0];
  GEN_28 = {1{$random}};
  req_typ = GEN_28[2:0];
  GEN_29 = {1{$random}};
  req_phys = GEN_29[0:0];
  GEN_30 = {2{$random}};
  req_data = GEN_30[63:0];
  GEN_31 = {2{$random}};
  grant_word = GEN_31[63:0];
  GEN_32 = {1{$random}};
  state = GEN_32[2:0];
  GEN_33 = {2{$random}};
  GEN_19 = GEN_33[63:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_1899) begin
        req_addr <= io_req_bits_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1899) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1899) begin
        req_cmd <= io_req_bits_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1899) begin
        req_typ <= io_req_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1899) begin
        req_phys <= io_req_bits_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1899) begin
        req_data <= io_req_bits_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1902) begin
        if(T_1762) begin
          grant_word <= T_1915;
        end
      end
    end
    if(reset) begin
      state <= 3'h0;
    end else begin
      if(T_1918) begin
        state <= 3'h0;
      end else begin
        if(T_1917) begin
          state <= 3'h4;
        end else begin
          if(T_1902) begin
            state <= 3'h3;
          end else begin
            if(T_1900) begin
              state <= 3'h2;
            end else begin
              if(T_1899) begin
                state <= 3'h1;
              end
            end
          end
        end
      end
    end
  end
endmodule
module MSHRFile(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [39:0] io_req_bits_addr,
  input  [8:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [63:0] io_req_bits_data,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  input   io_resp_ready,
  output  io_resp_valid,
  output [39:0] io_resp_bits_addr,
  output [8:0] io_resp_bits_tag,
  output [4:0] io_resp_bits_cmd,
  output [2:0] io_resp_bits_typ,
  output [63:0] io_resp_bits_data,
  output  io_resp_bits_replay,
  output  io_resp_bits_has_data,
  output [63:0] io_resp_bits_data_word_bypass,
  output [63:0] io_resp_bits_store_data,
  output  io_secondary_miss,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [11:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [8:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [63:0] io_replay_bits_data,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy,
  output  io_fence_rdy,
  output  io_replay_next
);
  wire [39:0] GEN_17;
  wire  T_2615;
  wire [39:0] GEN_18;
  wire  T_2617;
  wire  T_2618;
  reg [16:0] sdq_val;
  reg [31:0] GEN_5;
  wire [16:0] T_2622;
  wire  T_2623;
  wire  T_2624;
  wire  T_2625;
  wire  T_2626;
  wire  T_2627;
  wire  T_2628;
  wire  T_2629;
  wire  T_2630;
  wire  T_2631;
  wire  T_2632;
  wire  T_2633;
  wire  T_2634;
  wire  T_2635;
  wire  T_2636;
  wire  T_2637;
  wire  T_2638;
  wire  T_2639;
  wire [4:0] T_2657;
  wire [4:0] T_2658;
  wire [4:0] T_2659;
  wire [4:0] T_2660;
  wire [4:0] T_2661;
  wire [4:0] T_2662;
  wire [4:0] T_2663;
  wire [4:0] T_2664;
  wire [4:0] T_2665;
  wire [4:0] T_2666;
  wire [4:0] T_2667;
  wire [4:0] T_2668;
  wire [4:0] T_2669;
  wire [4:0] T_2670;
  wire [4:0] T_2671;
  wire [4:0] sdq_alloc_id;
  wire [16:0] GEN_19;
  wire  T_2674;
  wire  sdq_rdy;
  wire  T_2676;
  wire  T_2677;
  wire  T_2678;
  wire  T_2679;
  wire  T_2680;
  wire  T_2681;
  wire  T_2682;
  wire  T_2683;
  wire  T_2684;
  wire  sdq_enq;
  reg [63:0] sdq [0:16];
  reg [63:0] GEN_6;
  wire [63:0] sdq_T_4081_data;
  wire [4:0] sdq_T_4081_addr;
  wire  sdq_T_4081_en;
  wire [63:0] sdq_T_2686_data;
  wire [4:0] sdq_T_2686_addr;
  wire  sdq_T_2686_mask;
  wire  sdq_T_2686_en;
  wire  idxMatch_0;
  wire  idxMatch_1;
  wire [19:0] tagList_0;
  wire [19:0] tagList_1;
  wire [19:0] T_2702;
  wire [19:0] T_2704;
  wire [19:0] T_2706;
  wire [19:0] T_2707;
  wire [27:0] T_2708;
  wire [27:0] GEN_20;
  wire  tag_match;
  wire [19:0] wbTagList_0;
  wire [19:0] wbTagList_1;
  wire [3:0] refillMux_0_way_en;
  wire [11:0] refillMux_0_addr;
  wire [3:0] refillMux_1_way_en;
  wire [11:0] refillMux_1_addr;
  wire  meta_read_arb_clk;
  wire  meta_read_arb_reset;
  wire  meta_read_arb_io_in_0_ready;
  wire  meta_read_arb_io_in_0_valid;
  wire [5:0] meta_read_arb_io_in_0_bits_idx;
  wire [3:0] meta_read_arb_io_in_0_bits_way_en;
  wire [19:0] meta_read_arb_io_in_0_bits_tag;
  wire  meta_read_arb_io_in_1_ready;
  wire  meta_read_arb_io_in_1_valid;
  wire [5:0] meta_read_arb_io_in_1_bits_idx;
  wire [3:0] meta_read_arb_io_in_1_bits_way_en;
  wire [19:0] meta_read_arb_io_in_1_bits_tag;
  wire  meta_read_arb_io_out_ready;
  wire  meta_read_arb_io_out_valid;
  wire [5:0] meta_read_arb_io_out_bits_idx;
  wire [3:0] meta_read_arb_io_out_bits_way_en;
  wire [19:0] meta_read_arb_io_out_bits_tag;
  wire  meta_read_arb_io_chosen;
  wire  meta_write_arb_clk;
  wire  meta_write_arb_reset;
  wire  meta_write_arb_io_in_0_ready;
  wire  meta_write_arb_io_in_0_valid;
  wire [5:0] meta_write_arb_io_in_0_bits_idx;
  wire [3:0] meta_write_arb_io_in_0_bits_way_en;
  wire [19:0] meta_write_arb_io_in_0_bits_data_tag;
  wire [1:0] meta_write_arb_io_in_0_bits_data_coh_state;
  wire  meta_write_arb_io_in_1_ready;
  wire  meta_write_arb_io_in_1_valid;
  wire [5:0] meta_write_arb_io_in_1_bits_idx;
  wire [3:0] meta_write_arb_io_in_1_bits_way_en;
  wire [19:0] meta_write_arb_io_in_1_bits_data_tag;
  wire [1:0] meta_write_arb_io_in_1_bits_data_coh_state;
  wire  meta_write_arb_io_out_ready;
  wire  meta_write_arb_io_out_valid;
  wire [5:0] meta_write_arb_io_out_bits_idx;
  wire [3:0] meta_write_arb_io_out_bits_way_en;
  wire [19:0] meta_write_arb_io_out_bits_data_tag;
  wire [1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire  meta_write_arb_io_chosen;
  wire  mem_req_arb_clk;
  wire  mem_req_arb_reset;
  wire  mem_req_arb_io_in_0_ready;
  wire  mem_req_arb_io_in_0_valid;
  wire [25:0] mem_req_arb_io_in_0_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_0_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_0_bits_addr_beat;
  wire  mem_req_arb_io_in_0_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_0_bits_a_type;
  wire [11:0] mem_req_arb_io_in_0_bits_union;
  wire [63:0] mem_req_arb_io_in_0_bits_data;
  wire  mem_req_arb_io_in_1_ready;
  wire  mem_req_arb_io_in_1_valid;
  wire [25:0] mem_req_arb_io_in_1_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_1_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_1_bits_addr_beat;
  wire  mem_req_arb_io_in_1_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_1_bits_a_type;
  wire [11:0] mem_req_arb_io_in_1_bits_union;
  wire [63:0] mem_req_arb_io_in_1_bits_data;
  wire  mem_req_arb_io_in_2_ready;
  wire  mem_req_arb_io_in_2_valid;
  wire [25:0] mem_req_arb_io_in_2_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_2_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_2_bits_addr_beat;
  wire  mem_req_arb_io_in_2_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_2_bits_a_type;
  wire [11:0] mem_req_arb_io_in_2_bits_union;
  wire [63:0] mem_req_arb_io_in_2_bits_data;
  wire  mem_req_arb_io_out_ready;
  wire  mem_req_arb_io_out_valid;
  wire [25:0] mem_req_arb_io_out_bits_addr_block;
  wire [1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_out_bits_addr_beat;
  wire  mem_req_arb_io_out_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_out_bits_a_type;
  wire [11:0] mem_req_arb_io_out_bits_union;
  wire [63:0] mem_req_arb_io_out_bits_data;
  wire [1:0] mem_req_arb_io_chosen;
  wire  mem_finish_arb_clk;
  wire  mem_finish_arb_reset;
  wire  mem_finish_arb_io_in_0_ready;
  wire  mem_finish_arb_io_in_0_valid;
  wire [2:0] mem_finish_arb_io_in_0_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_0_bits_manager_id;
  wire  mem_finish_arb_io_in_1_ready;
  wire  mem_finish_arb_io_in_1_valid;
  wire [2:0] mem_finish_arb_io_in_1_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_1_bits_manager_id;
  wire  mem_finish_arb_io_in_2_ready;
  wire  mem_finish_arb_io_in_2_valid;
  wire [2:0] mem_finish_arb_io_in_2_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_2_bits_manager_id;
  wire  mem_finish_arb_io_out_ready;
  wire  mem_finish_arb_io_out_valid;
  wire [2:0] mem_finish_arb_io_out_bits_manager_xact_id;
  wire  mem_finish_arb_io_out_bits_manager_id;
  wire [1:0] mem_finish_arb_io_chosen;
  wire  wb_req_arb_clk;
  wire  wb_req_arb_reset;
  wire  wb_req_arb_io_in_0_ready;
  wire  wb_req_arb_io_in_0_valid;
  wire [2:0] wb_req_arb_io_in_0_bits_addr_beat;
  wire [25:0] wb_req_arb_io_in_0_bits_addr_block;
  wire [1:0] wb_req_arb_io_in_0_bits_client_xact_id;
  wire  wb_req_arb_io_in_0_bits_voluntary;
  wire [2:0] wb_req_arb_io_in_0_bits_r_type;
  wire [63:0] wb_req_arb_io_in_0_bits_data;
  wire [3:0] wb_req_arb_io_in_0_bits_way_en;
  wire  wb_req_arb_io_in_1_ready;
  wire  wb_req_arb_io_in_1_valid;
  wire [2:0] wb_req_arb_io_in_1_bits_addr_beat;
  wire [25:0] wb_req_arb_io_in_1_bits_addr_block;
  wire [1:0] wb_req_arb_io_in_1_bits_client_xact_id;
  wire  wb_req_arb_io_in_1_bits_voluntary;
  wire [2:0] wb_req_arb_io_in_1_bits_r_type;
  wire [63:0] wb_req_arb_io_in_1_bits_data;
  wire [3:0] wb_req_arb_io_in_1_bits_way_en;
  wire  wb_req_arb_io_out_ready;
  wire  wb_req_arb_io_out_valid;
  wire [2:0] wb_req_arb_io_out_bits_addr_beat;
  wire [25:0] wb_req_arb_io_out_bits_addr_block;
  wire [1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire  wb_req_arb_io_out_bits_voluntary;
  wire [2:0] wb_req_arb_io_out_bits_r_type;
  wire [63:0] wb_req_arb_io_out_bits_data;
  wire [3:0] wb_req_arb_io_out_bits_way_en;
  wire  wb_req_arb_io_chosen;
  wire  replay_arb_clk;
  wire  replay_arb_reset;
  wire  replay_arb_io_in_0_ready;
  wire  replay_arb_io_in_0_valid;
  wire [39:0] replay_arb_io_in_0_bits_addr;
  wire [8:0] replay_arb_io_in_0_bits_tag;
  wire [4:0] replay_arb_io_in_0_bits_cmd;
  wire [2:0] replay_arb_io_in_0_bits_typ;
  wire  replay_arb_io_in_0_bits_phys;
  wire [4:0] replay_arb_io_in_0_bits_sdq_id;
  wire  replay_arb_io_in_1_ready;
  wire  replay_arb_io_in_1_valid;
  wire [39:0] replay_arb_io_in_1_bits_addr;
  wire [8:0] replay_arb_io_in_1_bits_tag;
  wire [4:0] replay_arb_io_in_1_bits_cmd;
  wire [2:0] replay_arb_io_in_1_bits_typ;
  wire  replay_arb_io_in_1_bits_phys;
  wire [4:0] replay_arb_io_in_1_bits_sdq_id;
  wire  replay_arb_io_out_ready;
  wire  replay_arb_io_out_valid;
  wire [39:0] replay_arb_io_out_bits_addr;
  wire [8:0] replay_arb_io_out_bits_tag;
  wire [4:0] replay_arb_io_out_bits_cmd;
  wire [2:0] replay_arb_io_out_bits_typ;
  wire  replay_arb_io_out_bits_phys;
  wire [4:0] replay_arb_io_out_bits_sdq_id;
  wire  replay_arb_io_chosen;
  wire  alloc_arb_clk;
  wire  alloc_arb_reset;
  wire  alloc_arb_io_in_0_ready;
  wire  alloc_arb_io_in_0_valid;
  wire  alloc_arb_io_in_0_bits;
  wire  alloc_arb_io_in_1_ready;
  wire  alloc_arb_io_in_1_valid;
  wire  alloc_arb_io_in_1_bits;
  wire  alloc_arb_io_out_ready;
  wire  alloc_arb_io_out_valid;
  wire  alloc_arb_io_out_bits;
  wire  alloc_arb_io_chosen;
  wire  MSHR_2_clk;
  wire  MSHR_2_reset;
  wire  MSHR_2_io_req_pri_val;
  wire  MSHR_2_io_req_pri_rdy;
  wire  MSHR_2_io_req_sec_val;
  wire  MSHR_2_io_req_sec_rdy;
  wire [39:0] MSHR_2_io_req_bits_addr;
  wire [8:0] MSHR_2_io_req_bits_tag;
  wire [4:0] MSHR_2_io_req_bits_cmd;
  wire [2:0] MSHR_2_io_req_bits_typ;
  wire  MSHR_2_io_req_bits_phys;
  wire [4:0] MSHR_2_io_req_bits_sdq_id;
  wire  MSHR_2_io_req_bits_tag_match;
  wire [19:0] MSHR_2_io_req_bits_old_meta_tag;
  wire [1:0] MSHR_2_io_req_bits_old_meta_coh_state;
  wire [3:0] MSHR_2_io_req_bits_way_en;
  wire  MSHR_2_io_idx_match;
  wire [19:0] MSHR_2_io_tag;
  wire  MSHR_2_io_mem_req_ready;
  wire  MSHR_2_io_mem_req_valid;
  wire [25:0] MSHR_2_io_mem_req_bits_addr_block;
  wire [1:0] MSHR_2_io_mem_req_bits_client_xact_id;
  wire [2:0] MSHR_2_io_mem_req_bits_addr_beat;
  wire  MSHR_2_io_mem_req_bits_is_builtin_type;
  wire [2:0] MSHR_2_io_mem_req_bits_a_type;
  wire [11:0] MSHR_2_io_mem_req_bits_union;
  wire [63:0] MSHR_2_io_mem_req_bits_data;
  wire [3:0] MSHR_2_io_refill_way_en;
  wire [11:0] MSHR_2_io_refill_addr;
  wire  MSHR_2_io_meta_read_ready;
  wire  MSHR_2_io_meta_read_valid;
  wire [5:0] MSHR_2_io_meta_read_bits_idx;
  wire [3:0] MSHR_2_io_meta_read_bits_way_en;
  wire [19:0] MSHR_2_io_meta_read_bits_tag;
  wire  MSHR_2_io_meta_write_ready;
  wire  MSHR_2_io_meta_write_valid;
  wire [5:0] MSHR_2_io_meta_write_bits_idx;
  wire [3:0] MSHR_2_io_meta_write_bits_way_en;
  wire [19:0] MSHR_2_io_meta_write_bits_data_tag;
  wire [1:0] MSHR_2_io_meta_write_bits_data_coh_state;
  wire  MSHR_2_io_replay_ready;
  wire  MSHR_2_io_replay_valid;
  wire [39:0] MSHR_2_io_replay_bits_addr;
  wire [8:0] MSHR_2_io_replay_bits_tag;
  wire [4:0] MSHR_2_io_replay_bits_cmd;
  wire [2:0] MSHR_2_io_replay_bits_typ;
  wire  MSHR_2_io_replay_bits_phys;
  wire [4:0] MSHR_2_io_replay_bits_sdq_id;
  wire  MSHR_2_io_mem_grant_valid;
  wire [2:0] MSHR_2_io_mem_grant_bits_addr_beat;
  wire [1:0] MSHR_2_io_mem_grant_bits_client_xact_id;
  wire [2:0] MSHR_2_io_mem_grant_bits_manager_xact_id;
  wire  MSHR_2_io_mem_grant_bits_is_builtin_type;
  wire [3:0] MSHR_2_io_mem_grant_bits_g_type;
  wire [63:0] MSHR_2_io_mem_grant_bits_data;
  wire  MSHR_2_io_mem_grant_bits_manager_id;
  wire  MSHR_2_io_mem_finish_ready;
  wire  MSHR_2_io_mem_finish_valid;
  wire [2:0] MSHR_2_io_mem_finish_bits_manager_xact_id;
  wire  MSHR_2_io_mem_finish_bits_manager_id;
  wire  MSHR_2_io_wb_req_ready;
  wire  MSHR_2_io_wb_req_valid;
  wire [2:0] MSHR_2_io_wb_req_bits_addr_beat;
  wire [25:0] MSHR_2_io_wb_req_bits_addr_block;
  wire [1:0] MSHR_2_io_wb_req_bits_client_xact_id;
  wire  MSHR_2_io_wb_req_bits_voluntary;
  wire [2:0] MSHR_2_io_wb_req_bits_r_type;
  wire [63:0] MSHR_2_io_wb_req_bits_data;
  wire [3:0] MSHR_2_io_wb_req_bits_way_en;
  wire  MSHR_2_io_probe_rdy;
  wire [19:0] T_3871;
  wire  T_3872;
  wire  T_3873;
  wire [1:0] GEN_21;
  wire  T_3875;
  wire  T_3876;
  wire  T_3877;
  wire  T_3878;
  wire  T_3879;
  wire  T_3881;
  wire  GEN_7;
  wire  T_3884;
  wire  GEN_8;
  wire  MSHR_1_1_clk;
  wire  MSHR_1_1_reset;
  wire  MSHR_1_1_io_req_pri_val;
  wire  MSHR_1_1_io_req_pri_rdy;
  wire  MSHR_1_1_io_req_sec_val;
  wire  MSHR_1_1_io_req_sec_rdy;
  wire [39:0] MSHR_1_1_io_req_bits_addr;
  wire [8:0] MSHR_1_1_io_req_bits_tag;
  wire [4:0] MSHR_1_1_io_req_bits_cmd;
  wire [2:0] MSHR_1_1_io_req_bits_typ;
  wire  MSHR_1_1_io_req_bits_phys;
  wire [4:0] MSHR_1_1_io_req_bits_sdq_id;
  wire  MSHR_1_1_io_req_bits_tag_match;
  wire [19:0] MSHR_1_1_io_req_bits_old_meta_tag;
  wire [1:0] MSHR_1_1_io_req_bits_old_meta_coh_state;
  wire [3:0] MSHR_1_1_io_req_bits_way_en;
  wire  MSHR_1_1_io_idx_match;
  wire [19:0] MSHR_1_1_io_tag;
  wire  MSHR_1_1_io_mem_req_ready;
  wire  MSHR_1_1_io_mem_req_valid;
  wire [25:0] MSHR_1_1_io_mem_req_bits_addr_block;
  wire [1:0] MSHR_1_1_io_mem_req_bits_client_xact_id;
  wire [2:0] MSHR_1_1_io_mem_req_bits_addr_beat;
  wire  MSHR_1_1_io_mem_req_bits_is_builtin_type;
  wire [2:0] MSHR_1_1_io_mem_req_bits_a_type;
  wire [11:0] MSHR_1_1_io_mem_req_bits_union;
  wire [63:0] MSHR_1_1_io_mem_req_bits_data;
  wire [3:0] MSHR_1_1_io_refill_way_en;
  wire [11:0] MSHR_1_1_io_refill_addr;
  wire  MSHR_1_1_io_meta_read_ready;
  wire  MSHR_1_1_io_meta_read_valid;
  wire [5:0] MSHR_1_1_io_meta_read_bits_idx;
  wire [3:0] MSHR_1_1_io_meta_read_bits_way_en;
  wire [19:0] MSHR_1_1_io_meta_read_bits_tag;
  wire  MSHR_1_1_io_meta_write_ready;
  wire  MSHR_1_1_io_meta_write_valid;
  wire [5:0] MSHR_1_1_io_meta_write_bits_idx;
  wire [3:0] MSHR_1_1_io_meta_write_bits_way_en;
  wire [19:0] MSHR_1_1_io_meta_write_bits_data_tag;
  wire [1:0] MSHR_1_1_io_meta_write_bits_data_coh_state;
  wire  MSHR_1_1_io_replay_ready;
  wire  MSHR_1_1_io_replay_valid;
  wire [39:0] MSHR_1_1_io_replay_bits_addr;
  wire [8:0] MSHR_1_1_io_replay_bits_tag;
  wire [4:0] MSHR_1_1_io_replay_bits_cmd;
  wire [2:0] MSHR_1_1_io_replay_bits_typ;
  wire  MSHR_1_1_io_replay_bits_phys;
  wire [4:0] MSHR_1_1_io_replay_bits_sdq_id;
  wire  MSHR_1_1_io_mem_grant_valid;
  wire [2:0] MSHR_1_1_io_mem_grant_bits_addr_beat;
  wire [1:0] MSHR_1_1_io_mem_grant_bits_client_xact_id;
  wire [2:0] MSHR_1_1_io_mem_grant_bits_manager_xact_id;
  wire  MSHR_1_1_io_mem_grant_bits_is_builtin_type;
  wire [3:0] MSHR_1_1_io_mem_grant_bits_g_type;
  wire [63:0] MSHR_1_1_io_mem_grant_bits_data;
  wire  MSHR_1_1_io_mem_grant_bits_manager_id;
  wire  MSHR_1_1_io_mem_finish_ready;
  wire  MSHR_1_1_io_mem_finish_valid;
  wire [2:0] MSHR_1_1_io_mem_finish_bits_manager_xact_id;
  wire  MSHR_1_1_io_mem_finish_bits_manager_id;
  wire  MSHR_1_1_io_wb_req_ready;
  wire  MSHR_1_1_io_wb_req_valid;
  wire [2:0] MSHR_1_1_io_wb_req_bits_addr_beat;
  wire [25:0] MSHR_1_1_io_wb_req_bits_addr_block;
  wire [1:0] MSHR_1_1_io_wb_req_bits_client_xact_id;
  wire  MSHR_1_1_io_wb_req_bits_voluntary;
  wire [2:0] MSHR_1_1_io_wb_req_bits_r_type;
  wire [63:0] MSHR_1_1_io_wb_req_bits_data;
  wire [3:0] MSHR_1_1_io_wb_req_bits_way_en;
  wire  MSHR_1_1_io_probe_rdy;
  wire [19:0] T_3886;
  wire [1:0] GEN_22;
  wire  T_3890;
  wire  T_3891;
  wire  pri_rdy;
  wire  sec_rdy;
  wire  idx_match;
  wire  T_3893;
  wire  GEN_9;
  wire  T_3896;
  wire  GEN_10;
  wire  T_3899;
  wire  T_3901;
  wire  T_3902;
  wire  mmio_alloc_arb_clk;
  wire  mmio_alloc_arb_reset;
  wire  mmio_alloc_arb_io_in_0_ready;
  wire  mmio_alloc_arb_io_in_0_valid;
  wire  mmio_alloc_arb_io_in_0_bits;
  wire  mmio_alloc_arb_io_out_ready;
  wire  mmio_alloc_arb_io_out_valid;
  wire  mmio_alloc_arb_io_out_bits;
  wire  mmio_alloc_arb_io_chosen;
  wire  resp_arb_clk;
  wire  resp_arb_reset;
  wire  resp_arb_io_in_0_ready;
  wire  resp_arb_io_in_0_valid;
  wire [39:0] resp_arb_io_in_0_bits_addr;
  wire [8:0] resp_arb_io_in_0_bits_tag;
  wire [4:0] resp_arb_io_in_0_bits_cmd;
  wire [2:0] resp_arb_io_in_0_bits_typ;
  wire [63:0] resp_arb_io_in_0_bits_data;
  wire  resp_arb_io_in_0_bits_replay;
  wire  resp_arb_io_in_0_bits_has_data;
  wire [63:0] resp_arb_io_in_0_bits_data_word_bypass;
  wire [63:0] resp_arb_io_in_0_bits_store_data;
  wire  resp_arb_io_out_ready;
  wire  resp_arb_io_out_valid;
  wire [39:0] resp_arb_io_out_bits_addr;
  wire [8:0] resp_arb_io_out_bits_tag;
  wire [4:0] resp_arb_io_out_bits_cmd;
  wire [2:0] resp_arb_io_out_bits_typ;
  wire [63:0] resp_arb_io_out_bits_data;
  wire  resp_arb_io_out_bits_replay;
  wire  resp_arb_io_out_bits_has_data;
  wire [63:0] resp_arb_io_out_bits_data_word_bypass;
  wire [63:0] resp_arb_io_out_bits_store_data;
  wire  resp_arb_io_chosen;
  wire  IOMSHR_1_clk;
  wire  IOMSHR_1_reset;
  wire  IOMSHR_1_io_req_ready;
  wire  IOMSHR_1_io_req_valid;
  wire [39:0] IOMSHR_1_io_req_bits_addr;
  wire [8:0] IOMSHR_1_io_req_bits_tag;
  wire [4:0] IOMSHR_1_io_req_bits_cmd;
  wire [2:0] IOMSHR_1_io_req_bits_typ;
  wire  IOMSHR_1_io_req_bits_phys;
  wire [63:0] IOMSHR_1_io_req_bits_data;
  wire  IOMSHR_1_io_acquire_ready;
  wire  IOMSHR_1_io_acquire_valid;
  wire [25:0] IOMSHR_1_io_acquire_bits_addr_block;
  wire [1:0] IOMSHR_1_io_acquire_bits_client_xact_id;
  wire [2:0] IOMSHR_1_io_acquire_bits_addr_beat;
  wire  IOMSHR_1_io_acquire_bits_is_builtin_type;
  wire [2:0] IOMSHR_1_io_acquire_bits_a_type;
  wire [11:0] IOMSHR_1_io_acquire_bits_union;
  wire [63:0] IOMSHR_1_io_acquire_bits_data;
  wire  IOMSHR_1_io_grant_valid;
  wire [2:0] IOMSHR_1_io_grant_bits_addr_beat;
  wire [1:0] IOMSHR_1_io_grant_bits_client_xact_id;
  wire [2:0] IOMSHR_1_io_grant_bits_manager_xact_id;
  wire  IOMSHR_1_io_grant_bits_is_builtin_type;
  wire [3:0] IOMSHR_1_io_grant_bits_g_type;
  wire [63:0] IOMSHR_1_io_grant_bits_data;
  wire  IOMSHR_1_io_grant_bits_manager_id;
  wire  IOMSHR_1_io_finish_ready;
  wire  IOMSHR_1_io_finish_valid;
  wire [2:0] IOMSHR_1_io_finish_bits_manager_xact_id;
  wire  IOMSHR_1_io_finish_bits_manager_id;
  wire  IOMSHR_1_io_resp_ready;
  wire  IOMSHR_1_io_resp_valid;
  wire [39:0] IOMSHR_1_io_resp_bits_addr;
  wire [8:0] IOMSHR_1_io_resp_bits_tag;
  wire [4:0] IOMSHR_1_io_resp_bits_cmd;
  wire [2:0] IOMSHR_1_io_resp_bits_typ;
  wire [63:0] IOMSHR_1_io_resp_bits_data;
  wire  IOMSHR_1_io_resp_bits_replay;
  wire  IOMSHR_1_io_resp_bits_has_data;
  wire [63:0] IOMSHR_1_io_resp_bits_data_word_bypass;
  wire [63:0] IOMSHR_1_io_resp_bits_store_data;
  wire  IOMSHR_1_io_replay_next;
  wire  mmio_rdy;
  wire  T_3986;
  wire  T_3987;
  wire  T_3989;
  wire  GEN_11;
  wire  GEN_12;
  wire  T_3993;
  wire  T_3994;
  wire  T_3997;
  wire  T_3998;
  wire  T_3999;
  wire  T_4000;
  wire [3:0] GEN_0;
  wire [3:0] GEN_13;
  wire [11:0] GEN_1;
  wire [11:0] GEN_14;
  wire  T_4072;
  wire  T_4073;
  wire  T_4074;
  wire  T_4075;
  wire  T_4076;
  wire  T_4077;
  wire  T_4078;
  wire  T_4079;
  wire  free_sdq;
  reg [4:0] T_4080;
  reg [31:0] GEN_23;
  wire [4:0] GEN_15;
  wire  T_4082;
  wire [31:0] GEN_25;
  wire [31:0] T_4084;
  wire [16:0] GEN_26;
  wire [17:0] T_4086;
  wire [16:0] T_4087;
  wire [31:0] GEN_27;
  wire [31:0] T_4088;
  wire [31:0] T_4089;
  wire [31:0] GEN_28;
  wire [31:0] T_4090;
  wire [16:0] T_4129;
  wire [16:0] T_4130;
  wire [16:0] T_4131;
  wire [16:0] T_4132;
  wire [16:0] T_4133;
  wire [16:0] T_4134;
  wire [16:0] T_4135;
  wire [16:0] T_4136;
  wire [16:0] T_4137;
  wire [16:0] T_4138;
  wire [16:0] T_4139;
  wire [16:0] T_4140;
  wire [16:0] T_4141;
  wire [16:0] T_4142;
  wire [16:0] T_4143;
  wire [16:0] T_4144;
  wire [16:0] T_4145;
  wire [16:0] GEN_29;
  wire [17:0] T_4147;
  wire [16:0] T_4148;
  wire [16:0] T_4149;
  wire [31:0] GEN_30;
  wire [31:0] T_4150;
  wire [31:0] GEN_16;
  reg  GEN_2;
  reg [31:0] GEN_24;
  reg  GEN_3;
  reg [31:0] GEN_31;
  reg  GEN_4;
  reg [31:0] GEN_32;
  Arbiter meta_read_arb (
    .clk(meta_read_arb_clk),
    .reset(meta_read_arb_reset),
    .io_in_0_ready(meta_read_arb_io_in_0_ready),
    .io_in_0_valid(meta_read_arb_io_in_0_valid),
    .io_in_0_bits_idx(meta_read_arb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(meta_read_arb_io_in_0_bits_way_en),
    .io_in_0_bits_tag(meta_read_arb_io_in_0_bits_tag),
    .io_in_1_ready(meta_read_arb_io_in_1_ready),
    .io_in_1_valid(meta_read_arb_io_in_1_valid),
    .io_in_1_bits_idx(meta_read_arb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(meta_read_arb_io_in_1_bits_way_en),
    .io_in_1_bits_tag(meta_read_arb_io_in_1_bits_tag),
    .io_out_ready(meta_read_arb_io_out_ready),
    .io_out_valid(meta_read_arb_io_out_valid),
    .io_out_bits_idx(meta_read_arb_io_out_bits_idx),
    .io_out_bits_way_en(meta_read_arb_io_out_bits_way_en),
    .io_out_bits_tag(meta_read_arb_io_out_bits_tag),
    .io_chosen(meta_read_arb_io_chosen)
  );
  Arbiter_1 meta_write_arb (
    .clk(meta_write_arb_clk),
    .reset(meta_write_arb_reset),
    .io_in_0_ready(meta_write_arb_io_in_0_ready),
    .io_in_0_valid(meta_write_arb_io_in_0_valid),
    .io_in_0_bits_idx(meta_write_arb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(meta_write_arb_io_in_0_bits_way_en),
    .io_in_0_bits_data_tag(meta_write_arb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_coh_state(meta_write_arb_io_in_0_bits_data_coh_state),
    .io_in_1_ready(meta_write_arb_io_in_1_ready),
    .io_in_1_valid(meta_write_arb_io_in_1_valid),
    .io_in_1_bits_idx(meta_write_arb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(meta_write_arb_io_in_1_bits_way_en),
    .io_in_1_bits_data_tag(meta_write_arb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_coh_state(meta_write_arb_io_in_1_bits_data_coh_state),
    .io_out_ready(meta_write_arb_io_out_ready),
    .io_out_valid(meta_write_arb_io_out_valid),
    .io_out_bits_idx(meta_write_arb_io_out_bits_idx),
    .io_out_bits_way_en(meta_write_arb_io_out_bits_way_en),
    .io_out_bits_data_tag(meta_write_arb_io_out_bits_data_tag),
    .io_out_bits_data_coh_state(meta_write_arb_io_out_bits_data_coh_state),
    .io_chosen(meta_write_arb_io_chosen)
  );
  LockingArbiter mem_req_arb (
    .clk(mem_req_arb_clk),
    .reset(mem_req_arb_reset),
    .io_in_0_ready(mem_req_arb_io_in_0_ready),
    .io_in_0_valid(mem_req_arb_io_in_0_valid),
    .io_in_0_bits_addr_block(mem_req_arb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(mem_req_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(mem_req_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(mem_req_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(mem_req_arb_io_in_0_bits_a_type),
    .io_in_0_bits_union(mem_req_arb_io_in_0_bits_union),
    .io_in_0_bits_data(mem_req_arb_io_in_0_bits_data),
    .io_in_1_ready(mem_req_arb_io_in_1_ready),
    .io_in_1_valid(mem_req_arb_io_in_1_valid),
    .io_in_1_bits_addr_block(mem_req_arb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(mem_req_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(mem_req_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(mem_req_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(mem_req_arb_io_in_1_bits_a_type),
    .io_in_1_bits_union(mem_req_arb_io_in_1_bits_union),
    .io_in_1_bits_data(mem_req_arb_io_in_1_bits_data),
    .io_in_2_ready(mem_req_arb_io_in_2_ready),
    .io_in_2_valid(mem_req_arb_io_in_2_valid),
    .io_in_2_bits_addr_block(mem_req_arb_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(mem_req_arb_io_in_2_bits_client_xact_id),
    .io_in_2_bits_addr_beat(mem_req_arb_io_in_2_bits_addr_beat),
    .io_in_2_bits_is_builtin_type(mem_req_arb_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_a_type(mem_req_arb_io_in_2_bits_a_type),
    .io_in_2_bits_union(mem_req_arb_io_in_2_bits_union),
    .io_in_2_bits_data(mem_req_arb_io_in_2_bits_data),
    .io_out_ready(mem_req_arb_io_out_ready),
    .io_out_valid(mem_req_arb_io_out_valid),
    .io_out_bits_addr_block(mem_req_arb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(mem_req_arb_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(mem_req_arb_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(mem_req_arb_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(mem_req_arb_io_out_bits_a_type),
    .io_out_bits_union(mem_req_arb_io_out_bits_union),
    .io_out_bits_data(mem_req_arb_io_out_bits_data),
    .io_chosen(mem_req_arb_io_chosen)
  );
  Arbiter_2 mem_finish_arb (
    .clk(mem_finish_arb_clk),
    .reset(mem_finish_arb_reset),
    .io_in_0_ready(mem_finish_arb_io_in_0_ready),
    .io_in_0_valid(mem_finish_arb_io_in_0_valid),
    .io_in_0_bits_manager_xact_id(mem_finish_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_manager_id(mem_finish_arb_io_in_0_bits_manager_id),
    .io_in_1_ready(mem_finish_arb_io_in_1_ready),
    .io_in_1_valid(mem_finish_arb_io_in_1_valid),
    .io_in_1_bits_manager_xact_id(mem_finish_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_manager_id(mem_finish_arb_io_in_1_bits_manager_id),
    .io_in_2_ready(mem_finish_arb_io_in_2_ready),
    .io_in_2_valid(mem_finish_arb_io_in_2_valid),
    .io_in_2_bits_manager_xact_id(mem_finish_arb_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_manager_id(mem_finish_arb_io_in_2_bits_manager_id),
    .io_out_ready(mem_finish_arb_io_out_ready),
    .io_out_valid(mem_finish_arb_io_out_valid),
    .io_out_bits_manager_xact_id(mem_finish_arb_io_out_bits_manager_xact_id),
    .io_out_bits_manager_id(mem_finish_arb_io_out_bits_manager_id),
    .io_chosen(mem_finish_arb_io_chosen)
  );
  Arbiter_3 wb_req_arb (
    .clk(wb_req_arb_clk),
    .reset(wb_req_arb_reset),
    .io_in_0_ready(wb_req_arb_io_in_0_ready),
    .io_in_0_valid(wb_req_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(wb_req_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(wb_req_arb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(wb_req_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(wb_req_arb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(wb_req_arb_io_in_0_bits_r_type),
    .io_in_0_bits_data(wb_req_arb_io_in_0_bits_data),
    .io_in_0_bits_way_en(wb_req_arb_io_in_0_bits_way_en),
    .io_in_1_ready(wb_req_arb_io_in_1_ready),
    .io_in_1_valid(wb_req_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(wb_req_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(wb_req_arb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(wb_req_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(wb_req_arb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(wb_req_arb_io_in_1_bits_r_type),
    .io_in_1_bits_data(wb_req_arb_io_in_1_bits_data),
    .io_in_1_bits_way_en(wb_req_arb_io_in_1_bits_way_en),
    .io_out_ready(wb_req_arb_io_out_ready),
    .io_out_valid(wb_req_arb_io_out_valid),
    .io_out_bits_addr_beat(wb_req_arb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(wb_req_arb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(wb_req_arb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(wb_req_arb_io_out_bits_voluntary),
    .io_out_bits_r_type(wb_req_arb_io_out_bits_r_type),
    .io_out_bits_data(wb_req_arb_io_out_bits_data),
    .io_out_bits_way_en(wb_req_arb_io_out_bits_way_en),
    .io_chosen(wb_req_arb_io_chosen)
  );
  Arbiter_4 replay_arb (
    .clk(replay_arb_clk),
    .reset(replay_arb_reset),
    .io_in_0_ready(replay_arb_io_in_0_ready),
    .io_in_0_valid(replay_arb_io_in_0_valid),
    .io_in_0_bits_addr(replay_arb_io_in_0_bits_addr),
    .io_in_0_bits_tag(replay_arb_io_in_0_bits_tag),
    .io_in_0_bits_cmd(replay_arb_io_in_0_bits_cmd),
    .io_in_0_bits_typ(replay_arb_io_in_0_bits_typ),
    .io_in_0_bits_phys(replay_arb_io_in_0_bits_phys),
    .io_in_0_bits_sdq_id(replay_arb_io_in_0_bits_sdq_id),
    .io_in_1_ready(replay_arb_io_in_1_ready),
    .io_in_1_valid(replay_arb_io_in_1_valid),
    .io_in_1_bits_addr(replay_arb_io_in_1_bits_addr),
    .io_in_1_bits_tag(replay_arb_io_in_1_bits_tag),
    .io_in_1_bits_cmd(replay_arb_io_in_1_bits_cmd),
    .io_in_1_bits_typ(replay_arb_io_in_1_bits_typ),
    .io_in_1_bits_phys(replay_arb_io_in_1_bits_phys),
    .io_in_1_bits_sdq_id(replay_arb_io_in_1_bits_sdq_id),
    .io_out_ready(replay_arb_io_out_ready),
    .io_out_valid(replay_arb_io_out_valid),
    .io_out_bits_addr(replay_arb_io_out_bits_addr),
    .io_out_bits_tag(replay_arb_io_out_bits_tag),
    .io_out_bits_cmd(replay_arb_io_out_bits_cmd),
    .io_out_bits_typ(replay_arb_io_out_bits_typ),
    .io_out_bits_phys(replay_arb_io_out_bits_phys),
    .io_out_bits_sdq_id(replay_arb_io_out_bits_sdq_id),
    .io_chosen(replay_arb_io_chosen)
  );
  Arbiter_5 alloc_arb (
    .clk(alloc_arb_clk),
    .reset(alloc_arb_reset),
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_0_bits(alloc_arb_io_in_0_bits),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_in_1_bits(alloc_arb_io_in_1_bits),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid),
    .io_out_bits(alloc_arb_io_out_bits),
    .io_chosen(alloc_arb_io_chosen)
  );
  MSHR MSHR_2 (
    .clk(MSHR_2_clk),
    .reset(MSHR_2_reset),
    .io_req_pri_val(MSHR_2_io_req_pri_val),
    .io_req_pri_rdy(MSHR_2_io_req_pri_rdy),
    .io_req_sec_val(MSHR_2_io_req_sec_val),
    .io_req_sec_rdy(MSHR_2_io_req_sec_rdy),
    .io_req_bits_addr(MSHR_2_io_req_bits_addr),
    .io_req_bits_tag(MSHR_2_io_req_bits_tag),
    .io_req_bits_cmd(MSHR_2_io_req_bits_cmd),
    .io_req_bits_typ(MSHR_2_io_req_bits_typ),
    .io_req_bits_phys(MSHR_2_io_req_bits_phys),
    .io_req_bits_sdq_id(MSHR_2_io_req_bits_sdq_id),
    .io_req_bits_tag_match(MSHR_2_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(MSHR_2_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(MSHR_2_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(MSHR_2_io_req_bits_way_en),
    .io_idx_match(MSHR_2_io_idx_match),
    .io_tag(MSHR_2_io_tag),
    .io_mem_req_ready(MSHR_2_io_mem_req_ready),
    .io_mem_req_valid(MSHR_2_io_mem_req_valid),
    .io_mem_req_bits_addr_block(MSHR_2_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(MSHR_2_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(MSHR_2_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(MSHR_2_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(MSHR_2_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(MSHR_2_io_mem_req_bits_union),
    .io_mem_req_bits_data(MSHR_2_io_mem_req_bits_data),
    .io_refill_way_en(MSHR_2_io_refill_way_en),
    .io_refill_addr(MSHR_2_io_refill_addr),
    .io_meta_read_ready(MSHR_2_io_meta_read_ready),
    .io_meta_read_valid(MSHR_2_io_meta_read_valid),
    .io_meta_read_bits_idx(MSHR_2_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(MSHR_2_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(MSHR_2_io_meta_read_bits_tag),
    .io_meta_write_ready(MSHR_2_io_meta_write_ready),
    .io_meta_write_valid(MSHR_2_io_meta_write_valid),
    .io_meta_write_bits_idx(MSHR_2_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(MSHR_2_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(MSHR_2_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(MSHR_2_io_meta_write_bits_data_coh_state),
    .io_replay_ready(MSHR_2_io_replay_ready),
    .io_replay_valid(MSHR_2_io_replay_valid),
    .io_replay_bits_addr(MSHR_2_io_replay_bits_addr),
    .io_replay_bits_tag(MSHR_2_io_replay_bits_tag),
    .io_replay_bits_cmd(MSHR_2_io_replay_bits_cmd),
    .io_replay_bits_typ(MSHR_2_io_replay_bits_typ),
    .io_replay_bits_phys(MSHR_2_io_replay_bits_phys),
    .io_replay_bits_sdq_id(MSHR_2_io_replay_bits_sdq_id),
    .io_mem_grant_valid(MSHR_2_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(MSHR_2_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(MSHR_2_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(MSHR_2_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(MSHR_2_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(MSHR_2_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(MSHR_2_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(MSHR_2_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(MSHR_2_io_mem_finish_ready),
    .io_mem_finish_valid(MSHR_2_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(MSHR_2_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(MSHR_2_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(MSHR_2_io_wb_req_ready),
    .io_wb_req_valid(MSHR_2_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(MSHR_2_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(MSHR_2_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(MSHR_2_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(MSHR_2_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(MSHR_2_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(MSHR_2_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(MSHR_2_io_wb_req_bits_way_en),
    .io_probe_rdy(MSHR_2_io_probe_rdy)
  );
  MSHR_1 MSHR_1_1 (
    .clk(MSHR_1_1_clk),
    .reset(MSHR_1_1_reset),
    .io_req_pri_val(MSHR_1_1_io_req_pri_val),
    .io_req_pri_rdy(MSHR_1_1_io_req_pri_rdy),
    .io_req_sec_val(MSHR_1_1_io_req_sec_val),
    .io_req_sec_rdy(MSHR_1_1_io_req_sec_rdy),
    .io_req_bits_addr(MSHR_1_1_io_req_bits_addr),
    .io_req_bits_tag(MSHR_1_1_io_req_bits_tag),
    .io_req_bits_cmd(MSHR_1_1_io_req_bits_cmd),
    .io_req_bits_typ(MSHR_1_1_io_req_bits_typ),
    .io_req_bits_phys(MSHR_1_1_io_req_bits_phys),
    .io_req_bits_sdq_id(MSHR_1_1_io_req_bits_sdq_id),
    .io_req_bits_tag_match(MSHR_1_1_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(MSHR_1_1_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(MSHR_1_1_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(MSHR_1_1_io_req_bits_way_en),
    .io_idx_match(MSHR_1_1_io_idx_match),
    .io_tag(MSHR_1_1_io_tag),
    .io_mem_req_ready(MSHR_1_1_io_mem_req_ready),
    .io_mem_req_valid(MSHR_1_1_io_mem_req_valid),
    .io_mem_req_bits_addr_block(MSHR_1_1_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(MSHR_1_1_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(MSHR_1_1_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(MSHR_1_1_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(MSHR_1_1_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(MSHR_1_1_io_mem_req_bits_union),
    .io_mem_req_bits_data(MSHR_1_1_io_mem_req_bits_data),
    .io_refill_way_en(MSHR_1_1_io_refill_way_en),
    .io_refill_addr(MSHR_1_1_io_refill_addr),
    .io_meta_read_ready(MSHR_1_1_io_meta_read_ready),
    .io_meta_read_valid(MSHR_1_1_io_meta_read_valid),
    .io_meta_read_bits_idx(MSHR_1_1_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(MSHR_1_1_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(MSHR_1_1_io_meta_read_bits_tag),
    .io_meta_write_ready(MSHR_1_1_io_meta_write_ready),
    .io_meta_write_valid(MSHR_1_1_io_meta_write_valid),
    .io_meta_write_bits_idx(MSHR_1_1_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(MSHR_1_1_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(MSHR_1_1_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(MSHR_1_1_io_meta_write_bits_data_coh_state),
    .io_replay_ready(MSHR_1_1_io_replay_ready),
    .io_replay_valid(MSHR_1_1_io_replay_valid),
    .io_replay_bits_addr(MSHR_1_1_io_replay_bits_addr),
    .io_replay_bits_tag(MSHR_1_1_io_replay_bits_tag),
    .io_replay_bits_cmd(MSHR_1_1_io_replay_bits_cmd),
    .io_replay_bits_typ(MSHR_1_1_io_replay_bits_typ),
    .io_replay_bits_phys(MSHR_1_1_io_replay_bits_phys),
    .io_replay_bits_sdq_id(MSHR_1_1_io_replay_bits_sdq_id),
    .io_mem_grant_valid(MSHR_1_1_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(MSHR_1_1_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(MSHR_1_1_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(MSHR_1_1_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(MSHR_1_1_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(MSHR_1_1_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(MSHR_1_1_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(MSHR_1_1_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(MSHR_1_1_io_mem_finish_ready),
    .io_mem_finish_valid(MSHR_1_1_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(MSHR_1_1_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(MSHR_1_1_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(MSHR_1_1_io_wb_req_ready),
    .io_wb_req_valid(MSHR_1_1_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(MSHR_1_1_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(MSHR_1_1_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(MSHR_1_1_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(MSHR_1_1_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(MSHR_1_1_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(MSHR_1_1_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(MSHR_1_1_io_wb_req_bits_way_en),
    .io_probe_rdy(MSHR_1_1_io_probe_rdy)
  );
  Arbiter_6 mmio_alloc_arb (
    .clk(mmio_alloc_arb_clk),
    .reset(mmio_alloc_arb_reset),
    .io_in_0_ready(mmio_alloc_arb_io_in_0_ready),
    .io_in_0_valid(mmio_alloc_arb_io_in_0_valid),
    .io_in_0_bits(mmio_alloc_arb_io_in_0_bits),
    .io_out_ready(mmio_alloc_arb_io_out_ready),
    .io_out_valid(mmio_alloc_arb_io_out_valid),
    .io_out_bits(mmio_alloc_arb_io_out_bits),
    .io_chosen(mmio_alloc_arb_io_chosen)
  );
  Arbiter_7 resp_arb (
    .clk(resp_arb_clk),
    .reset(resp_arb_reset),
    .io_in_0_ready(resp_arb_io_in_0_ready),
    .io_in_0_valid(resp_arb_io_in_0_valid),
    .io_in_0_bits_addr(resp_arb_io_in_0_bits_addr),
    .io_in_0_bits_tag(resp_arb_io_in_0_bits_tag),
    .io_in_0_bits_cmd(resp_arb_io_in_0_bits_cmd),
    .io_in_0_bits_typ(resp_arb_io_in_0_bits_typ),
    .io_in_0_bits_data(resp_arb_io_in_0_bits_data),
    .io_in_0_bits_replay(resp_arb_io_in_0_bits_replay),
    .io_in_0_bits_has_data(resp_arb_io_in_0_bits_has_data),
    .io_in_0_bits_data_word_bypass(resp_arb_io_in_0_bits_data_word_bypass),
    .io_in_0_bits_store_data(resp_arb_io_in_0_bits_store_data),
    .io_out_ready(resp_arb_io_out_ready),
    .io_out_valid(resp_arb_io_out_valid),
    .io_out_bits_addr(resp_arb_io_out_bits_addr),
    .io_out_bits_tag(resp_arb_io_out_bits_tag),
    .io_out_bits_cmd(resp_arb_io_out_bits_cmd),
    .io_out_bits_typ(resp_arb_io_out_bits_typ),
    .io_out_bits_data(resp_arb_io_out_bits_data),
    .io_out_bits_replay(resp_arb_io_out_bits_replay),
    .io_out_bits_has_data(resp_arb_io_out_bits_has_data),
    .io_out_bits_data_word_bypass(resp_arb_io_out_bits_data_word_bypass),
    .io_out_bits_store_data(resp_arb_io_out_bits_store_data),
    .io_chosen(resp_arb_io_chosen)
  );
  IOMSHR IOMSHR_1 (
    .clk(IOMSHR_1_clk),
    .reset(IOMSHR_1_reset),
    .io_req_ready(IOMSHR_1_io_req_ready),
    .io_req_valid(IOMSHR_1_io_req_valid),
    .io_req_bits_addr(IOMSHR_1_io_req_bits_addr),
    .io_req_bits_tag(IOMSHR_1_io_req_bits_tag),
    .io_req_bits_cmd(IOMSHR_1_io_req_bits_cmd),
    .io_req_bits_typ(IOMSHR_1_io_req_bits_typ),
    .io_req_bits_phys(IOMSHR_1_io_req_bits_phys),
    .io_req_bits_data(IOMSHR_1_io_req_bits_data),
    .io_acquire_ready(IOMSHR_1_io_acquire_ready),
    .io_acquire_valid(IOMSHR_1_io_acquire_valid),
    .io_acquire_bits_addr_block(IOMSHR_1_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(IOMSHR_1_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(IOMSHR_1_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(IOMSHR_1_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(IOMSHR_1_io_acquire_bits_a_type),
    .io_acquire_bits_union(IOMSHR_1_io_acquire_bits_union),
    .io_acquire_bits_data(IOMSHR_1_io_acquire_bits_data),
    .io_grant_valid(IOMSHR_1_io_grant_valid),
    .io_grant_bits_addr_beat(IOMSHR_1_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(IOMSHR_1_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(IOMSHR_1_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(IOMSHR_1_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(IOMSHR_1_io_grant_bits_g_type),
    .io_grant_bits_data(IOMSHR_1_io_grant_bits_data),
    .io_grant_bits_manager_id(IOMSHR_1_io_grant_bits_manager_id),
    .io_finish_ready(IOMSHR_1_io_finish_ready),
    .io_finish_valid(IOMSHR_1_io_finish_valid),
    .io_finish_bits_manager_xact_id(IOMSHR_1_io_finish_bits_manager_xact_id),
    .io_finish_bits_manager_id(IOMSHR_1_io_finish_bits_manager_id),
    .io_resp_ready(IOMSHR_1_io_resp_ready),
    .io_resp_valid(IOMSHR_1_io_resp_valid),
    .io_resp_bits_addr(IOMSHR_1_io_resp_bits_addr),
    .io_resp_bits_tag(IOMSHR_1_io_resp_bits_tag),
    .io_resp_bits_cmd(IOMSHR_1_io_resp_bits_cmd),
    .io_resp_bits_typ(IOMSHR_1_io_resp_bits_typ),
    .io_resp_bits_data(IOMSHR_1_io_resp_bits_data),
    .io_resp_bits_replay(IOMSHR_1_io_resp_bits_replay),
    .io_resp_bits_has_data(IOMSHR_1_io_resp_bits_has_data),
    .io_resp_bits_data_word_bypass(IOMSHR_1_io_resp_bits_data_word_bypass),
    .io_resp_bits_store_data(IOMSHR_1_io_resp_bits_store_data),
    .io_replay_next(IOMSHR_1_io_replay_next)
  );
  assign io_req_ready = T_4000;
  assign io_resp_valid = resp_arb_io_out_valid;
  assign io_resp_bits_addr = resp_arb_io_out_bits_addr;
  assign io_resp_bits_tag = resp_arb_io_out_bits_tag;
  assign io_resp_bits_cmd = resp_arb_io_out_bits_cmd;
  assign io_resp_bits_typ = resp_arb_io_out_bits_typ;
  assign io_resp_bits_data = resp_arb_io_out_bits_data;
  assign io_resp_bits_replay = resp_arb_io_out_bits_replay;
  assign io_resp_bits_has_data = resp_arb_io_out_bits_has_data;
  assign io_resp_bits_data_word_bypass = resp_arb_io_out_bits_data_word_bypass;
  assign io_resp_bits_store_data = resp_arb_io_out_bits_store_data;
  assign io_secondary_miss = idx_match;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_mem_req_bits_addr_block = mem_req_arb_io_out_bits_addr_block;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr_beat = mem_req_arb_io_out_bits_addr_beat;
  assign io_mem_req_bits_is_builtin_type = mem_req_arb_io_out_bits_is_builtin_type;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_union = mem_req_arb_io_out_bits_union;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_refill_way_en = GEN_0;
  assign io_refill_addr = GEN_1;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_bits_way_en = meta_read_arb_io_out_bits_way_en;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_data = sdq_T_4081_data;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_mem_finish_bits_manager_xact_id = mem_finish_arb_io_out_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = mem_finish_arb_io_out_bits_manager_id;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_wb_req_bits_addr_beat = wb_req_arb_io_out_bits_addr_beat;
  assign io_wb_req_bits_addr_block = wb_req_arb_io_out_bits_addr_block;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_voluntary = wb_req_arb_io_out_bits_voluntary;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_data = wb_req_arb_io_out_bits_data;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_probe_rdy = GEN_10;
  assign io_fence_rdy = GEN_11;
  assign io_replay_next = GEN_12;
  assign GEN_17 = {{8'd0}, 32'h80000000};
  assign T_2615 = GEN_17 <= io_req_bits_addr;
  assign GEN_18 = {{7'd0}, 33'h100000000};
  assign T_2617 = io_req_bits_addr < GEN_18;
  assign T_2618 = T_2615 & T_2617;
  assign T_2622 = ~ sdq_val;
  assign T_2623 = T_2622[0];
  assign T_2624 = T_2622[1];
  assign T_2625 = T_2622[2];
  assign T_2626 = T_2622[3];
  assign T_2627 = T_2622[4];
  assign T_2628 = T_2622[5];
  assign T_2629 = T_2622[6];
  assign T_2630 = T_2622[7];
  assign T_2631 = T_2622[8];
  assign T_2632 = T_2622[9];
  assign T_2633 = T_2622[10];
  assign T_2634 = T_2622[11];
  assign T_2635 = T_2622[12];
  assign T_2636 = T_2622[13];
  assign T_2637 = T_2622[14];
  assign T_2638 = T_2622[15];
  assign T_2639 = T_2622[16];
  assign T_2657 = T_2638 ? {{1'd0}, 4'hf} : 5'h10;
  assign T_2658 = T_2637 ? {{1'd0}, 4'he} : T_2657;
  assign T_2659 = T_2636 ? {{1'd0}, 4'hd} : T_2658;
  assign T_2660 = T_2635 ? {{1'd0}, 4'hc} : T_2659;
  assign T_2661 = T_2634 ? {{1'd0}, 4'hb} : T_2660;
  assign T_2662 = T_2633 ? {{1'd0}, 4'ha} : T_2661;
  assign T_2663 = T_2632 ? {{1'd0}, 4'h9} : T_2662;
  assign T_2664 = T_2631 ? {{1'd0}, 4'h8} : T_2663;
  assign T_2665 = T_2630 ? {{2'd0}, 3'h7} : T_2664;
  assign T_2666 = T_2629 ? {{2'd0}, 3'h6} : T_2665;
  assign T_2667 = T_2628 ? {{2'd0}, 3'h5} : T_2666;
  assign T_2668 = T_2627 ? {{2'd0}, 3'h4} : T_2667;
  assign T_2669 = T_2626 ? {{3'd0}, 2'h3} : T_2668;
  assign T_2670 = T_2625 ? {{3'd0}, 2'h2} : T_2669;
  assign T_2671 = T_2624 ? {{4'd0}, 1'h1} : T_2670;
  assign sdq_alloc_id = T_2623 ? {{4'd0}, 1'h0} : T_2671;
  assign GEN_19 = {{16'd0}, 1'h0};
  assign T_2674 = T_2622 == GEN_19;
  assign sdq_rdy = T_2674 == 1'h0;
  assign T_2676 = io_req_valid & io_req_ready;
  assign T_2677 = T_2676 & T_2618;
  assign T_2678 = io_req_bits_cmd == 5'h1;
  assign T_2679 = io_req_bits_cmd == 5'h7;
  assign T_2680 = T_2678 | T_2679;
  assign T_2681 = io_req_bits_cmd[3];
  assign T_2682 = io_req_bits_cmd == 5'h4;
  assign T_2683 = T_2681 | T_2682;
  assign T_2684 = T_2680 | T_2683;
  assign sdq_enq = T_2677 & T_2684;
  assign sdq_T_4081_addr = T_4080;
  assign sdq_T_4081_en = 1'h1;
  `ifdef SYNTHESIS
  assign sdq_T_4081_data = sdq[sdq_T_4081_addr];
  `else
  assign sdq_T_4081_data = sdq_T_4081_addr >= 5'h11 ? $random : sdq[sdq_T_4081_addr];
  `endif
  assign sdq_T_2686_data = io_req_bits_data;
  assign sdq_T_2686_addr = sdq_alloc_id;
  assign sdq_T_2686_mask = sdq_enq;
  assign sdq_T_2686_en = sdq_enq;
  assign idxMatch_0 = MSHR_2_io_idx_match;
  assign idxMatch_1 = MSHR_1_1_io_idx_match;
  assign tagList_0 = MSHR_2_io_tag;
  assign tagList_1 = MSHR_1_1_io_tag;
  assign T_2702 = idxMatch_0 ? tagList_0 : {{19'd0}, 1'h0};
  assign T_2704 = idxMatch_1 ? tagList_1 : {{19'd0}, 1'h0};
  assign T_2706 = T_2702 | T_2704;
  assign T_2707 = T_2706;
  assign T_2708 = io_req_bits_addr[39:12];
  assign GEN_20 = {{8'd0}, T_2707};
  assign tag_match = GEN_20 == T_2708;
  assign wbTagList_0 = T_3871;
  assign wbTagList_1 = T_3886;
  assign refillMux_0_way_en = MSHR_2_io_refill_way_en;
  assign refillMux_0_addr = MSHR_2_io_refill_addr;
  assign refillMux_1_way_en = MSHR_1_1_io_refill_way_en;
  assign refillMux_1_addr = MSHR_1_1_io_refill_addr;
  assign meta_read_arb_clk = clk;
  assign meta_read_arb_reset = reset;
  assign meta_read_arb_io_in_0_valid = MSHR_2_io_meta_read_valid;
  assign meta_read_arb_io_in_0_bits_idx = MSHR_2_io_meta_read_bits_idx;
  assign meta_read_arb_io_in_0_bits_way_en = MSHR_2_io_meta_read_bits_way_en;
  assign meta_read_arb_io_in_0_bits_tag = MSHR_2_io_meta_read_bits_tag;
  assign meta_read_arb_io_in_1_valid = MSHR_1_1_io_meta_read_valid;
  assign meta_read_arb_io_in_1_bits_idx = MSHR_1_1_io_meta_read_bits_idx;
  assign meta_read_arb_io_in_1_bits_way_en = MSHR_1_1_io_meta_read_bits_way_en;
  assign meta_read_arb_io_in_1_bits_tag = MSHR_1_1_io_meta_read_bits_tag;
  assign meta_read_arb_io_out_ready = io_meta_read_ready;
  assign meta_write_arb_clk = clk;
  assign meta_write_arb_reset = reset;
  assign meta_write_arb_io_in_0_valid = MSHR_2_io_meta_write_valid;
  assign meta_write_arb_io_in_0_bits_idx = MSHR_2_io_meta_write_bits_idx;
  assign meta_write_arb_io_in_0_bits_way_en = MSHR_2_io_meta_write_bits_way_en;
  assign meta_write_arb_io_in_0_bits_data_tag = MSHR_2_io_meta_write_bits_data_tag;
  assign meta_write_arb_io_in_0_bits_data_coh_state = MSHR_2_io_meta_write_bits_data_coh_state;
  assign meta_write_arb_io_in_1_valid = MSHR_1_1_io_meta_write_valid;
  assign meta_write_arb_io_in_1_bits_idx = MSHR_1_1_io_meta_write_bits_idx;
  assign meta_write_arb_io_in_1_bits_way_en = MSHR_1_1_io_meta_write_bits_way_en;
  assign meta_write_arb_io_in_1_bits_data_tag = MSHR_1_1_io_meta_write_bits_data_tag;
  assign meta_write_arb_io_in_1_bits_data_coh_state = MSHR_1_1_io_meta_write_bits_data_coh_state;
  assign meta_write_arb_io_out_ready = io_meta_write_ready;
  assign mem_req_arb_clk = clk;
  assign mem_req_arb_reset = reset;
  assign mem_req_arb_io_in_0_valid = MSHR_2_io_mem_req_valid;
  assign mem_req_arb_io_in_0_bits_addr_block = MSHR_2_io_mem_req_bits_addr_block;
  assign mem_req_arb_io_in_0_bits_client_xact_id = MSHR_2_io_mem_req_bits_client_xact_id;
  assign mem_req_arb_io_in_0_bits_addr_beat = MSHR_2_io_mem_req_bits_addr_beat;
  assign mem_req_arb_io_in_0_bits_is_builtin_type = MSHR_2_io_mem_req_bits_is_builtin_type;
  assign mem_req_arb_io_in_0_bits_a_type = MSHR_2_io_mem_req_bits_a_type;
  assign mem_req_arb_io_in_0_bits_union = MSHR_2_io_mem_req_bits_union;
  assign mem_req_arb_io_in_0_bits_data = MSHR_2_io_mem_req_bits_data;
  assign mem_req_arb_io_in_1_valid = MSHR_1_1_io_mem_req_valid;
  assign mem_req_arb_io_in_1_bits_addr_block = MSHR_1_1_io_mem_req_bits_addr_block;
  assign mem_req_arb_io_in_1_bits_client_xact_id = MSHR_1_1_io_mem_req_bits_client_xact_id;
  assign mem_req_arb_io_in_1_bits_addr_beat = MSHR_1_1_io_mem_req_bits_addr_beat;
  assign mem_req_arb_io_in_1_bits_is_builtin_type = MSHR_1_1_io_mem_req_bits_is_builtin_type;
  assign mem_req_arb_io_in_1_bits_a_type = MSHR_1_1_io_mem_req_bits_a_type;
  assign mem_req_arb_io_in_1_bits_union = MSHR_1_1_io_mem_req_bits_union;
  assign mem_req_arb_io_in_1_bits_data = MSHR_1_1_io_mem_req_bits_data;
  assign mem_req_arb_io_in_2_valid = IOMSHR_1_io_acquire_valid;
  assign mem_req_arb_io_in_2_bits_addr_block = IOMSHR_1_io_acquire_bits_addr_block;
  assign mem_req_arb_io_in_2_bits_client_xact_id = IOMSHR_1_io_acquire_bits_client_xact_id;
  assign mem_req_arb_io_in_2_bits_addr_beat = IOMSHR_1_io_acquire_bits_addr_beat;
  assign mem_req_arb_io_in_2_bits_is_builtin_type = IOMSHR_1_io_acquire_bits_is_builtin_type;
  assign mem_req_arb_io_in_2_bits_a_type = IOMSHR_1_io_acquire_bits_a_type;
  assign mem_req_arb_io_in_2_bits_union = IOMSHR_1_io_acquire_bits_union;
  assign mem_req_arb_io_in_2_bits_data = IOMSHR_1_io_acquire_bits_data;
  assign mem_req_arb_io_out_ready = io_mem_req_ready;
  assign mem_finish_arb_clk = clk;
  assign mem_finish_arb_reset = reset;
  assign mem_finish_arb_io_in_0_valid = MSHR_2_io_mem_finish_valid;
  assign mem_finish_arb_io_in_0_bits_manager_xact_id = MSHR_2_io_mem_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_0_bits_manager_id = MSHR_2_io_mem_finish_bits_manager_id;
  assign mem_finish_arb_io_in_1_valid = MSHR_1_1_io_mem_finish_valid;
  assign mem_finish_arb_io_in_1_bits_manager_xact_id = MSHR_1_1_io_mem_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_1_bits_manager_id = MSHR_1_1_io_mem_finish_bits_manager_id;
  assign mem_finish_arb_io_in_2_valid = IOMSHR_1_io_finish_valid;
  assign mem_finish_arb_io_in_2_bits_manager_xact_id = IOMSHR_1_io_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_2_bits_manager_id = IOMSHR_1_io_finish_bits_manager_id;
  assign mem_finish_arb_io_out_ready = io_mem_finish_ready;
  assign wb_req_arb_clk = clk;
  assign wb_req_arb_reset = reset;
  assign wb_req_arb_io_in_0_valid = MSHR_2_io_wb_req_valid;
  assign wb_req_arb_io_in_0_bits_addr_beat = MSHR_2_io_wb_req_bits_addr_beat;
  assign wb_req_arb_io_in_0_bits_addr_block = MSHR_2_io_wb_req_bits_addr_block;
  assign wb_req_arb_io_in_0_bits_client_xact_id = MSHR_2_io_wb_req_bits_client_xact_id;
  assign wb_req_arb_io_in_0_bits_voluntary = MSHR_2_io_wb_req_bits_voluntary;
  assign wb_req_arb_io_in_0_bits_r_type = MSHR_2_io_wb_req_bits_r_type;
  assign wb_req_arb_io_in_0_bits_data = MSHR_2_io_wb_req_bits_data;
  assign wb_req_arb_io_in_0_bits_way_en = MSHR_2_io_wb_req_bits_way_en;
  assign wb_req_arb_io_in_1_valid = MSHR_1_1_io_wb_req_valid;
  assign wb_req_arb_io_in_1_bits_addr_beat = MSHR_1_1_io_wb_req_bits_addr_beat;
  assign wb_req_arb_io_in_1_bits_addr_block = MSHR_1_1_io_wb_req_bits_addr_block;
  assign wb_req_arb_io_in_1_bits_client_xact_id = MSHR_1_1_io_wb_req_bits_client_xact_id;
  assign wb_req_arb_io_in_1_bits_voluntary = MSHR_1_1_io_wb_req_bits_voluntary;
  assign wb_req_arb_io_in_1_bits_r_type = MSHR_1_1_io_wb_req_bits_r_type;
  assign wb_req_arb_io_in_1_bits_data = MSHR_1_1_io_wb_req_bits_data;
  assign wb_req_arb_io_in_1_bits_way_en = MSHR_1_1_io_wb_req_bits_way_en;
  assign wb_req_arb_io_out_ready = io_wb_req_ready;
  assign replay_arb_clk = clk;
  assign replay_arb_reset = reset;
  assign replay_arb_io_in_0_valid = MSHR_2_io_replay_valid;
  assign replay_arb_io_in_0_bits_addr = MSHR_2_io_replay_bits_addr;
  assign replay_arb_io_in_0_bits_tag = MSHR_2_io_replay_bits_tag;
  assign replay_arb_io_in_0_bits_cmd = MSHR_2_io_replay_bits_cmd;
  assign replay_arb_io_in_0_bits_typ = MSHR_2_io_replay_bits_typ;
  assign replay_arb_io_in_0_bits_phys = MSHR_2_io_replay_bits_phys;
  assign replay_arb_io_in_0_bits_sdq_id = MSHR_2_io_replay_bits_sdq_id;
  assign replay_arb_io_in_1_valid = MSHR_1_1_io_replay_valid;
  assign replay_arb_io_in_1_bits_addr = MSHR_1_1_io_replay_bits_addr;
  assign replay_arb_io_in_1_bits_tag = MSHR_1_1_io_replay_bits_tag;
  assign replay_arb_io_in_1_bits_cmd = MSHR_1_1_io_replay_bits_cmd;
  assign replay_arb_io_in_1_bits_typ = MSHR_1_1_io_replay_bits_typ;
  assign replay_arb_io_in_1_bits_phys = MSHR_1_1_io_replay_bits_phys;
  assign replay_arb_io_in_1_bits_sdq_id = MSHR_1_1_io_replay_bits_sdq_id;
  assign replay_arb_io_out_ready = io_replay_ready;
  assign alloc_arb_clk = clk;
  assign alloc_arb_reset = reset;
  assign alloc_arb_io_in_0_valid = MSHR_2_io_req_pri_rdy;
  assign alloc_arb_io_in_0_bits = GEN_2;
  assign alloc_arb_io_in_1_valid = MSHR_1_1_io_req_pri_rdy;
  assign alloc_arb_io_in_1_bits = GEN_3;
  assign alloc_arb_io_out_ready = T_3902;
  assign MSHR_2_clk = clk;
  assign MSHR_2_reset = reset;
  assign MSHR_2_io_req_pri_val = alloc_arb_io_in_0_ready;
  assign MSHR_2_io_req_sec_val = T_3873;
  assign MSHR_2_io_req_bits_addr = io_req_bits_addr;
  assign MSHR_2_io_req_bits_tag = io_req_bits_tag;
  assign MSHR_2_io_req_bits_cmd = io_req_bits_cmd;
  assign MSHR_2_io_req_bits_typ = io_req_bits_typ;
  assign MSHR_2_io_req_bits_phys = io_req_bits_phys;
  assign MSHR_2_io_req_bits_sdq_id = sdq_alloc_id;
  assign MSHR_2_io_req_bits_tag_match = io_req_bits_tag_match;
  assign MSHR_2_io_req_bits_old_meta_tag = io_req_bits_old_meta_tag;
  assign MSHR_2_io_req_bits_old_meta_coh_state = io_req_bits_old_meta_coh_state;
  assign MSHR_2_io_req_bits_way_en = io_req_bits_way_en;
  assign MSHR_2_io_mem_req_ready = mem_req_arb_io_in_0_ready;
  assign MSHR_2_io_meta_read_ready = meta_read_arb_io_in_0_ready;
  assign MSHR_2_io_meta_write_ready = meta_write_arb_io_in_0_ready;
  assign MSHR_2_io_replay_ready = replay_arb_io_in_0_ready;
  assign MSHR_2_io_mem_grant_valid = T_3876;
  assign MSHR_2_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign MSHR_2_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign MSHR_2_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign MSHR_2_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign MSHR_2_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign MSHR_2_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign MSHR_2_io_mem_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign MSHR_2_io_mem_finish_ready = mem_finish_arb_io_in_0_ready;
  assign MSHR_2_io_wb_req_ready = wb_req_arb_io_in_0_ready;
  assign T_3871 = MSHR_2_io_wb_req_bits_addr_block[25:6];
  assign T_3872 = io_req_valid & sdq_rdy;
  assign T_3873 = T_3872 & tag_match;
  assign GEN_21 = {{1'd0}, 1'h0};
  assign T_3875 = io_mem_grant_bits_client_xact_id == GEN_21;
  assign T_3876 = io_mem_grant_valid & T_3875;
  assign T_3877 = MSHR_2_io_req_pri_rdy;
  assign T_3878 = MSHR_2_io_req_sec_rdy;
  assign T_3879 = MSHR_2_io_idx_match;
  assign T_3881 = MSHR_2_io_req_pri_rdy == 1'h0;
  assign GEN_7 = T_3881 ? 1'h0 : 1'h1;
  assign T_3884 = MSHR_2_io_probe_rdy == 1'h0;
  assign GEN_8 = T_3884 ? 1'h0 : 1'h1;
  assign MSHR_1_1_clk = clk;
  assign MSHR_1_1_reset = reset;
  assign MSHR_1_1_io_req_pri_val = alloc_arb_io_in_1_ready;
  assign MSHR_1_1_io_req_sec_val = T_3873;
  assign MSHR_1_1_io_req_bits_addr = io_req_bits_addr;
  assign MSHR_1_1_io_req_bits_tag = io_req_bits_tag;
  assign MSHR_1_1_io_req_bits_cmd = io_req_bits_cmd;
  assign MSHR_1_1_io_req_bits_typ = io_req_bits_typ;
  assign MSHR_1_1_io_req_bits_phys = io_req_bits_phys;
  assign MSHR_1_1_io_req_bits_sdq_id = sdq_alloc_id;
  assign MSHR_1_1_io_req_bits_tag_match = io_req_bits_tag_match;
  assign MSHR_1_1_io_req_bits_old_meta_tag = io_req_bits_old_meta_tag;
  assign MSHR_1_1_io_req_bits_old_meta_coh_state = io_req_bits_old_meta_coh_state;
  assign MSHR_1_1_io_req_bits_way_en = io_req_bits_way_en;
  assign MSHR_1_1_io_mem_req_ready = mem_req_arb_io_in_1_ready;
  assign MSHR_1_1_io_meta_read_ready = meta_read_arb_io_in_1_ready;
  assign MSHR_1_1_io_meta_write_ready = meta_write_arb_io_in_1_ready;
  assign MSHR_1_1_io_replay_ready = replay_arb_io_in_1_ready;
  assign MSHR_1_1_io_mem_grant_valid = T_3891;
  assign MSHR_1_1_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign MSHR_1_1_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign MSHR_1_1_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign MSHR_1_1_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign MSHR_1_1_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign MSHR_1_1_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign MSHR_1_1_io_mem_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign MSHR_1_1_io_mem_finish_ready = mem_finish_arb_io_in_1_ready;
  assign MSHR_1_1_io_wb_req_ready = wb_req_arb_io_in_1_ready;
  assign T_3886 = MSHR_1_1_io_wb_req_bits_addr_block[25:6];
  assign GEN_22 = {{1'd0}, 1'h1};
  assign T_3890 = io_mem_grant_bits_client_xact_id == GEN_22;
  assign T_3891 = io_mem_grant_valid & T_3890;
  assign pri_rdy = T_3877 | MSHR_1_1_io_req_pri_rdy;
  assign sec_rdy = T_3878 | MSHR_1_1_io_req_sec_rdy;
  assign idx_match = T_3879 | MSHR_1_1_io_idx_match;
  assign T_3893 = MSHR_1_1_io_req_pri_rdy == 1'h0;
  assign GEN_9 = T_3893 ? 1'h0 : GEN_7;
  assign T_3896 = MSHR_1_1_io_probe_rdy == 1'h0;
  assign GEN_10 = T_3896 ? 1'h0 : GEN_8;
  assign T_3899 = T_3872 & T_2618;
  assign T_3901 = idx_match == 1'h0;
  assign T_3902 = T_3899 & T_3901;
  assign mmio_alloc_arb_clk = clk;
  assign mmio_alloc_arb_reset = reset;
  assign mmio_alloc_arb_io_in_0_valid = IOMSHR_1_io_req_ready;
  assign mmio_alloc_arb_io_in_0_bits = GEN_4;
  assign mmio_alloc_arb_io_out_ready = T_3994;
  assign resp_arb_clk = clk;
  assign resp_arb_reset = reset;
  assign resp_arb_io_in_0_valid = IOMSHR_1_io_resp_valid;
  assign resp_arb_io_in_0_bits_addr = IOMSHR_1_io_resp_bits_addr;
  assign resp_arb_io_in_0_bits_tag = IOMSHR_1_io_resp_bits_tag;
  assign resp_arb_io_in_0_bits_cmd = IOMSHR_1_io_resp_bits_cmd;
  assign resp_arb_io_in_0_bits_typ = IOMSHR_1_io_resp_bits_typ;
  assign resp_arb_io_in_0_bits_data = IOMSHR_1_io_resp_bits_data;
  assign resp_arb_io_in_0_bits_replay = IOMSHR_1_io_resp_bits_replay;
  assign resp_arb_io_in_0_bits_has_data = IOMSHR_1_io_resp_bits_has_data;
  assign resp_arb_io_in_0_bits_data_word_bypass = IOMSHR_1_io_resp_bits_data_word_bypass;
  assign resp_arb_io_in_0_bits_store_data = IOMSHR_1_io_resp_bits_store_data;
  assign resp_arb_io_out_ready = io_resp_ready;
  assign IOMSHR_1_clk = clk;
  assign IOMSHR_1_reset = reset;
  assign IOMSHR_1_io_req_valid = mmio_alloc_arb_io_in_0_ready;
  assign IOMSHR_1_io_req_bits_addr = io_req_bits_addr;
  assign IOMSHR_1_io_req_bits_tag = io_req_bits_tag;
  assign IOMSHR_1_io_req_bits_cmd = io_req_bits_cmd;
  assign IOMSHR_1_io_req_bits_typ = io_req_bits_typ;
  assign IOMSHR_1_io_req_bits_phys = io_req_bits_phys;
  assign IOMSHR_1_io_req_bits_data = io_req_bits_data;
  assign IOMSHR_1_io_acquire_ready = mem_req_arb_io_in_2_ready;
  assign IOMSHR_1_io_grant_valid = T_3987;
  assign IOMSHR_1_io_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign IOMSHR_1_io_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign IOMSHR_1_io_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign IOMSHR_1_io_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign IOMSHR_1_io_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign IOMSHR_1_io_grant_bits_data = io_mem_grant_bits_data;
  assign IOMSHR_1_io_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign IOMSHR_1_io_finish_ready = mem_finish_arb_io_in_2_ready;
  assign IOMSHR_1_io_resp_ready = resp_arb_io_in_0_ready;
  assign mmio_rdy = IOMSHR_1_io_req_ready;
  assign T_3986 = io_mem_grant_bits_client_xact_id == 2'h2;
  assign T_3987 = io_mem_grant_valid & T_3986;
  assign T_3989 = IOMSHR_1_io_req_ready == 1'h0;
  assign GEN_11 = T_3989 ? 1'h0 : GEN_9;
  assign GEN_12 = IOMSHR_1_io_replay_next;
  assign T_3993 = T_2618 == 1'h0;
  assign T_3994 = io_req_valid & T_3993;
  assign T_3997 = tag_match & sec_rdy;
  assign T_3998 = idx_match ? T_3997 : pri_rdy;
  assign T_3999 = T_3998 & sdq_rdy;
  assign T_4000 = T_3993 ? mmio_rdy : T_3999;
  assign GEN_0 = GEN_13;
  assign GEN_13 = GEN_22 == io_mem_grant_bits_client_xact_id ? refillMux_1_way_en : refillMux_0_way_en;
  assign GEN_1 = GEN_14;
  assign GEN_14 = GEN_22 == io_mem_grant_bits_client_xact_id ? refillMux_1_addr : refillMux_0_addr;
  assign T_4072 = io_replay_ready & io_replay_valid;
  assign T_4073 = io_replay_bits_cmd == 5'h1;
  assign T_4074 = io_replay_bits_cmd == 5'h7;
  assign T_4075 = T_4073 | T_4074;
  assign T_4076 = io_replay_bits_cmd[3];
  assign T_4077 = io_replay_bits_cmd == 5'h4;
  assign T_4078 = T_4076 | T_4077;
  assign T_4079 = T_4075 | T_4078;
  assign free_sdq = T_4072 & T_4079;
  assign GEN_15 = free_sdq ? replay_arb_io_out_bits_sdq_id : T_4080;
  assign T_4082 = io_replay_valid | sdq_enq;
  assign GEN_25 = {{31'd0}, 1'h1};
  assign T_4084 = GEN_25 << replay_arb_io_out_bits_sdq_id;
  assign GEN_26 = {{16'd0}, free_sdq};
  assign T_4086 = 17'h0 - GEN_26;
  assign T_4087 = T_4086[16:0];
  assign GEN_27 = {{15'd0}, T_4087};
  assign T_4088 = T_4084 & GEN_27;
  assign T_4089 = ~ T_4088;
  assign GEN_28 = {{15'd0}, sdq_val};
  assign T_4090 = GEN_28 & T_4089;
  assign T_4129 = T_2639 ? 17'h10000 : 17'h0;
  assign T_4130 = T_2638 ? 17'h8000 : T_4129;
  assign T_4131 = T_2637 ? 17'h4000 : T_4130;
  assign T_4132 = T_2636 ? 17'h2000 : T_4131;
  assign T_4133 = T_2635 ? 17'h1000 : T_4132;
  assign T_4134 = T_2634 ? 17'h800 : T_4133;
  assign T_4135 = T_2633 ? 17'h400 : T_4134;
  assign T_4136 = T_2632 ? 17'h200 : T_4135;
  assign T_4137 = T_2631 ? 17'h100 : T_4136;
  assign T_4138 = T_2630 ? 17'h80 : T_4137;
  assign T_4139 = T_2629 ? 17'h40 : T_4138;
  assign T_4140 = T_2628 ? 17'h20 : T_4139;
  assign T_4141 = T_2627 ? 17'h10 : T_4140;
  assign T_4142 = T_2626 ? 17'h8 : T_4141;
  assign T_4143 = T_2625 ? 17'h4 : T_4142;
  assign T_4144 = T_2624 ? 17'h2 : T_4143;
  assign T_4145 = T_2623 ? 17'h1 : T_4144;
  assign GEN_29 = {{16'd0}, sdq_enq};
  assign T_4147 = 17'h0 - GEN_29;
  assign T_4148 = T_4147[16:0];
  assign T_4149 = T_4145 & T_4148;
  assign GEN_30 = {{15'd0}, T_4149};
  assign T_4150 = T_4090 | GEN_30;
  assign GEN_16 = T_4082 ? T_4150 : {{15'd0}, sdq_val};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_5 = {1{$random}};
  sdq_val = GEN_5[16:0];
  GEN_6 = {2{$random}};
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    sdq[initvar] = GEN_6[63:0];
  GEN_23 = {1{$random}};
  T_4080 = GEN_23[4:0];
  GEN_24 = {1{$random}};
  GEN_2 = GEN_24[0:0];
  GEN_31 = {1{$random}};
  GEN_3 = GEN_31[0:0];
  GEN_32 = {1{$random}};
  GEN_4 = GEN_32[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      sdq_val <= 17'h0;
    end else begin
      sdq_val <= GEN_16[16:0];
    end
    if(sdq_T_2686_en & sdq_T_2686_mask) begin
      sdq[sdq_T_2686_addr] <= sdq_T_2686_data;
    end
    if(1'h0) begin
    end else begin
      if(free_sdq) begin
        T_4080 <= replay_arb_io_out_bits_sdq_id;
      end
    end
  end
endmodule
module MetadataArray(
  input   clk,
  input   reset,
  output  io_read_ready,
  input   io_read_valid,
  input  [5:0] io_read_bits_idx,
  input  [3:0] io_read_bits_way_en,
  output  io_write_ready,
  input   io_write_valid,
  input  [5:0] io_write_bits_idx,
  input  [3:0] io_write_bits_way_en,
  input  [19:0] io_write_bits_data_tag,
  input  [1:0] io_write_bits_data_coh_state,
  output [19:0] io_resp_0_tag,
  output [1:0] io_resp_0_coh_state,
  output [19:0] io_resp_1_tag,
  output [1:0] io_resp_1_coh_state,
  output [19:0] io_resp_2_tag,
  output [1:0] io_resp_2_coh_state,
  output [19:0] io_resp_3_tag,
  output [1:0] io_resp_3_coh_state
);
  wire [1:0] T_50_state;
  wire [19:0] rstVal_tag;
  wire [1:0] rstVal_coh_state;
  reg [6:0] rst_cnt;
  reg [31:0] GEN_1;
  wire  rst;
  wire [6:0] waddr;
  wire [19:0] T_2358_tag;
  wire [1:0] T_2358_coh_state;
  wire [21:0] wdata;
  wire [3:0] T_2457;
  wire  GEN_25;
  wire [3:0] T_2458;
  wire  T_2459;
  wire  T_2460;
  wire  T_2461;
  wire  T_2462;
  wire [6:0] GEN_27;
  wire [7:0] T_2473;
  wire [6:0] T_2474;
  wire [6:0] GEN_0;
  reg [21:0] T_2483_0 [0:63];
  reg [31:0] GEN_2;
  wire [21:0] T_2483_0_T_2500_data;
  wire [5:0] T_2483_0_T_2500_addr;
  wire  T_2483_0_T_2500_en;
  reg [5:0] GEN_3;
  reg [31:0] GEN_4;
  reg  GEN_5;
  reg [31:0] GEN_6;
  wire [21:0] T_2483_0_T_2494_data;
  wire [5:0] T_2483_0_T_2494_addr;
  wire  T_2483_0_T_2494_mask;
  wire  T_2483_0_T_2494_en;
  reg [21:0] T_2483_1 [0:63];
  reg [31:0] GEN_7;
  wire [21:0] T_2483_1_T_2500_data;
  wire [5:0] T_2483_1_T_2500_addr;
  wire  T_2483_1_T_2500_en;
  reg [5:0] GEN_8;
  reg [31:0] GEN_9;
  reg  GEN_10;
  reg [31:0] GEN_11;
  wire [21:0] T_2483_1_T_2494_data;
  wire [5:0] T_2483_1_T_2494_addr;
  wire  T_2483_1_T_2494_mask;
  wire  T_2483_1_T_2494_en;
  reg [21:0] T_2483_2 [0:63];
  reg [31:0] GEN_12;
  wire [21:0] T_2483_2_T_2500_data;
  wire [5:0] T_2483_2_T_2500_addr;
  wire  T_2483_2_T_2500_en;
  reg [5:0] GEN_13;
  reg [31:0] GEN_14;
  reg  GEN_15;
  reg [31:0] GEN_16;
  wire [21:0] T_2483_2_T_2494_data;
  wire [5:0] T_2483_2_T_2494_addr;
  wire  T_2483_2_T_2494_mask;
  wire  T_2483_2_T_2494_en;
  reg [21:0] T_2483_3 [0:63];
  reg [31:0] GEN_18;
  wire [21:0] T_2483_3_T_2500_data;
  wire [5:0] T_2483_3_T_2500_addr;
  wire  T_2483_3_T_2500_en;
  reg [5:0] GEN_20;
  reg [31:0] GEN_22;
  reg  GEN_24;
  reg [31:0] GEN_26;
  wire [21:0] T_2483_3_T_2494_data;
  wire [5:0] T_2483_3_T_2494_addr;
  wire  T_2483_3_T_2494_mask;
  wire  T_2483_3_T_2494_en;
  wire  T_2484;
  wire [21:0] T_2490_0;
  wire [21:0] T_2490_1;
  wire [21:0] T_2490_2;
  wire [21:0] T_2490_3;
  wire  GEN_17;
  wire  GEN_19;
  wire  GEN_21;
  wire  GEN_23;
  wire [5:0] T_2497;
  wire [43:0] T_2502;
  wire [43:0] T_2503;
  wire [87:0] T_2504;
  wire [19:0] T_3366_0_tag;
  wire [1:0] T_3366_0_coh_state;
  wire [19:0] T_3366_1_tag;
  wire [1:0] T_3366_1_coh_state;
  wire [19:0] T_3366_2_tag;
  wire [1:0] T_3366_2_coh_state;
  wire [19:0] T_3366_3_tag;
  wire [1:0] T_3366_3_coh_state;
  wire [1:0] T_3843;
  wire [19:0] T_3844;
  wire [1:0] T_3845;
  wire [19:0] T_3846;
  wire [1:0] T_3847;
  wire [19:0] T_3848;
  wire [1:0] T_3849;
  wire [19:0] T_3850;
  wire  T_3852;
  wire  T_3854;
  wire  T_3855;
  assign io_read_ready = T_3855;
  assign io_write_ready = T_3852;
  assign io_resp_0_tag = T_3366_0_tag;
  assign io_resp_0_coh_state = T_3366_0_coh_state;
  assign io_resp_1_tag = T_3366_1_tag;
  assign io_resp_1_coh_state = T_3366_1_coh_state;
  assign io_resp_2_tag = T_3366_2_tag;
  assign io_resp_2_coh_state = T_3366_2_coh_state;
  assign io_resp_3_tag = T_3366_3_tag;
  assign io_resp_3_coh_state = T_3366_3_coh_state;
  assign T_50_state = {{1'd0}, 1'h0};
  assign rstVal_tag = {{19'd0}, 1'h0};
  assign rstVal_coh_state = T_50_state;
  assign rst = rst_cnt < 7'h40;
  assign waddr = rst ? rst_cnt : {{1'd0}, io_write_bits_idx};
  assign T_2358_tag = rst ? rstVal_tag : io_write_bits_data_tag;
  assign T_2358_coh_state = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign wdata = {T_2358_tag,T_2358_coh_state};
  assign T_2457 = $signed(io_write_bits_way_en);
  assign GEN_25 = $signed(1'h1);
  assign T_2458 = rst ? $signed({4{GEN_25}}) : $signed(T_2457);
  assign T_2459 = T_2458[0];
  assign T_2460 = T_2458[1];
  assign T_2461 = T_2458[2];
  assign T_2462 = T_2458[3];
  assign GEN_27 = {{6'd0}, 1'h1};
  assign T_2473 = rst_cnt + GEN_27;
  assign T_2474 = T_2473[6:0];
  assign GEN_0 = rst ? T_2474 : rst_cnt;
  assign T_2483_0_T_2500_addr = T_2497;
  assign T_2483_0_T_2500_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_2483_0_T_2500_data = T_2483_0[GEN_3];
  `else
  assign T_2483_0_T_2500_data = GEN_3 >= 7'h40 ? $random : T_2483_0[GEN_3];
  `endif
  assign T_2483_0_T_2494_data = T_2490_0;
  assign T_2483_0_T_2494_addr = waddr[5:0];
  assign T_2483_0_T_2494_mask = GEN_17;
  assign T_2483_0_T_2494_en = T_2484;
  assign T_2483_1_T_2500_addr = T_2497;
  assign T_2483_1_T_2500_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_2483_1_T_2500_data = T_2483_1[GEN_8];
  `else
  assign T_2483_1_T_2500_data = GEN_8 >= 7'h40 ? $random : T_2483_1[GEN_8];
  `endif
  assign T_2483_1_T_2494_data = T_2490_1;
  assign T_2483_1_T_2494_addr = waddr[5:0];
  assign T_2483_1_T_2494_mask = GEN_19;
  assign T_2483_1_T_2494_en = T_2484;
  assign T_2483_2_T_2500_addr = T_2497;
  assign T_2483_2_T_2500_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_2483_2_T_2500_data = T_2483_2[GEN_13];
  `else
  assign T_2483_2_T_2500_data = GEN_13 >= 7'h40 ? $random : T_2483_2[GEN_13];
  `endif
  assign T_2483_2_T_2494_data = T_2490_2;
  assign T_2483_2_T_2494_addr = waddr[5:0];
  assign T_2483_2_T_2494_mask = GEN_21;
  assign T_2483_2_T_2494_en = T_2484;
  assign T_2483_3_T_2500_addr = T_2497;
  assign T_2483_3_T_2500_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_2483_3_T_2500_data = T_2483_3[GEN_20];
  `else
  assign T_2483_3_T_2500_data = GEN_20 >= 7'h40 ? $random : T_2483_3[GEN_20];
  `endif
  assign T_2483_3_T_2494_data = T_2490_3;
  assign T_2483_3_T_2494_addr = waddr[5:0];
  assign T_2483_3_T_2494_mask = GEN_23;
  assign T_2483_3_T_2494_en = T_2484;
  assign T_2484 = rst | io_write_valid;
  assign T_2490_0 = wdata;
  assign T_2490_1 = wdata;
  assign T_2490_2 = wdata;
  assign T_2490_3 = wdata;
  assign GEN_17 = T_2484 ? T_2459 : 1'h0;
  assign GEN_19 = T_2484 ? T_2460 : 1'h0;
  assign GEN_21 = T_2484 ? T_2461 : 1'h0;
  assign GEN_23 = T_2484 ? T_2462 : 1'h0;
  assign T_2497 = io_read_bits_idx;
  assign T_2502 = {T_2483_1_T_2500_data,T_2483_0_T_2500_data};
  assign T_2503 = {T_2483_3_T_2500_data,T_2483_2_T_2500_data};
  assign T_2504 = {T_2503,T_2502};
  assign T_3366_0_tag = T_3844;
  assign T_3366_0_coh_state = T_3843;
  assign T_3366_1_tag = T_3846;
  assign T_3366_1_coh_state = T_3845;
  assign T_3366_2_tag = T_3848;
  assign T_3366_2_coh_state = T_3847;
  assign T_3366_3_tag = T_3850;
  assign T_3366_3_coh_state = T_3849;
  assign T_3843 = T_2504[1:0];
  assign T_3844 = T_2504[21:2];
  assign T_3845 = T_2504[23:22];
  assign T_3846 = T_2504[43:24];
  assign T_3847 = T_2504[45:44];
  assign T_3848 = T_2504[65:46];
  assign T_3849 = T_2504[67:66];
  assign T_3850 = T_2504[87:68];
  assign T_3852 = rst == 1'h0;
  assign T_3854 = io_write_valid == 1'h0;
  assign T_3855 = T_3852 & T_3854;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_1 = {1{$random}};
  rst_cnt = GEN_1[6:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2483_0[initvar] = GEN_2[21:0];
  GEN_4 = {1{$random}};
  GEN_3 = GEN_4[5:0];
  GEN_6 = {1{$random}};
  GEN_5 = GEN_6[0:0];
  GEN_7 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2483_1[initvar] = GEN_7[21:0];
  GEN_9 = {1{$random}};
  GEN_8 = GEN_9[5:0];
  GEN_11 = {1{$random}};
  GEN_10 = GEN_11[0:0];
  GEN_12 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2483_2[initvar] = GEN_12[21:0];
  GEN_14 = {1{$random}};
  GEN_13 = GEN_14[5:0];
  GEN_16 = {1{$random}};
  GEN_15 = GEN_16[0:0];
  GEN_18 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2483_3[initvar] = GEN_18[21:0];
  GEN_22 = {1{$random}};
  GEN_20 = GEN_22[5:0];
  GEN_26 = {1{$random}};
  GEN_24 = GEN_26[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else begin
      if(rst) begin
        rst_cnt <= T_2474;
      end
    end
    GEN_3 <= T_2483_0_T_2500_addr;
    GEN_5 <= T_2483_0_T_2500_en;
    if(T_2483_0_T_2494_en & T_2483_0_T_2494_mask) begin
      T_2483_0[T_2483_0_T_2494_addr] <= T_2483_0_T_2494_data;
    end
    GEN_8 <= T_2483_1_T_2500_addr;
    GEN_10 <= T_2483_1_T_2500_en;
    if(T_2483_1_T_2494_en & T_2483_1_T_2494_mask) begin
      T_2483_1[T_2483_1_T_2494_addr] <= T_2483_1_T_2494_data;
    end
    GEN_13 <= T_2483_2_T_2500_addr;
    GEN_15 <= T_2483_2_T_2500_en;
    if(T_2483_2_T_2494_en & T_2483_2_T_2494_mask) begin
      T_2483_2[T_2483_2_T_2494_addr] <= T_2483_2_T_2494_data;
    end
    GEN_20 <= T_2483_3_T_2500_addr;
    GEN_24 <= T_2483_3_T_2500_en;
    if(T_2483_3_T_2494_en & T_2483_3_T_2494_mask) begin
      T_2483_3[T_2483_3_T_2494_addr] <= T_2483_3_T_2494_data;
    end
  end
endmodule
module Arbiter_8(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [5:0] io_in_2_bits_idx,
  input  [3:0] io_in_2_bits_way_en,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [5:0] io_in_3_bits_idx,
  input  [3:0] io_in_3_bits_way_en,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [5:0] io_in_4_bits_idx,
  input  [3:0] io_in_4_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [2:0] io_chosen
);
  wire [2:0] GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [2:0] GEN_3;
  wire [5:0] GEN_4;
  wire [3:0] GEN_5;
  wire [2:0] GEN_6;
  wire [5:0] GEN_7;
  wire [3:0] GEN_8;
  wire [2:0] GEN_9;
  wire [5:0] GEN_10;
  wire [3:0] GEN_11;
  wire  T_934;
  wire  T_935;
  wire  T_936;
  wire  T_938;
  wire  T_940;
  wire  T_942;
  wire  T_944;
  wire  T_946;
  wire  T_947;
  wire  T_948;
  wire  T_949;
  wire  T_951;
  wire  T_952;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_946;
  assign io_in_2_ready = T_947;
  assign io_in_3_ready = T_948;
  assign io_in_4_ready = T_949;
  assign io_out_valid = T_952;
  assign io_out_bits_idx = GEN_10;
  assign io_out_bits_way_en = GEN_11;
  assign io_chosen = GEN_9;
  assign GEN_0 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_1 = io_in_3_valid ? io_in_3_bits_idx : io_in_4_bits_idx;
  assign GEN_2 = io_in_3_valid ? io_in_3_bits_way_en : io_in_4_bits_way_en;
  assign GEN_3 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_0;
  assign GEN_4 = io_in_2_valid ? io_in_2_bits_idx : GEN_1;
  assign GEN_5 = io_in_2_valid ? io_in_2_bits_way_en : GEN_2;
  assign GEN_6 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_3;
  assign GEN_7 = io_in_1_valid ? io_in_1_bits_idx : GEN_4;
  assign GEN_8 = io_in_1_valid ? io_in_1_bits_way_en : GEN_5;
  assign GEN_9 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_6;
  assign GEN_10 = io_in_0_valid ? io_in_0_bits_idx : GEN_7;
  assign GEN_11 = io_in_0_valid ? io_in_0_bits_way_en : GEN_8;
  assign T_934 = io_in_0_valid | io_in_1_valid;
  assign T_935 = T_934 | io_in_2_valid;
  assign T_936 = T_935 | io_in_3_valid;
  assign T_938 = io_in_0_valid == 1'h0;
  assign T_940 = T_934 == 1'h0;
  assign T_942 = T_935 == 1'h0;
  assign T_944 = T_936 == 1'h0;
  assign T_946 = T_938 & io_out_ready;
  assign T_947 = T_940 & io_out_ready;
  assign T_948 = T_942 & io_out_ready;
  assign T_949 = T_944 & io_out_ready;
  assign T_951 = T_944 == 1'h0;
  assign T_952 = T_951 | io_in_4_valid;
endmodule
module DataArray(
  input   clk,
  input   reset,
  output  io_read_ready,
  input   io_read_valid,
  input  [3:0] io_read_bits_way_en,
  input  [11:0] io_read_bits_addr,
  output  io_write_ready,
  input   io_write_valid,
  input  [3:0] io_write_bits_way_en,
  input  [11:0] io_write_bits_addr,
  input   io_write_bits_wmask,
  input  [63:0] io_write_bits_data,
  output [63:0] io_resp_0,
  output [63:0] io_resp_1,
  output [63:0] io_resp_2,
  output [63:0] io_resp_3
);
  wire [8:0] waddr;
  wire [8:0] raddr;
  wire  T_815;
  wire [63:0] T_823_0;
  reg [11:0] T_825;
  reg [31:0] GEN_1;
  wire [11:0] GEN_0;
  reg [63:0] T_834_0 [0:511];
  reg [63:0] GEN_2;
  wire [63:0] T_834_0_T_860_data;
  wire [8:0] T_834_0_T_860_addr;
  wire  T_834_0_T_860_en;
  reg [8:0] GEN_3;
  reg [31:0] GEN_4;
  reg  GEN_5;
  reg [31:0] GEN_6;
  wire [63:0] T_834_0_T_851_data;
  wire [8:0] T_834_0_T_851_addr;
  wire  T_834_0_T_851_mask;
  wire  T_834_0_T_851_en;
  wire  T_837;
  wire  T_839;
  wire [63:0] T_846_0;
  wire  GEN_8;
  wire [8:0] T_857;
  wire [63:0] T_868_0;
  wire  T_870;
  wire [63:0] T_878_0;
  reg [11:0] T_880;
  reg [31:0] GEN_7;
  wire [11:0] GEN_10;
  reg [63:0] T_889_0 [0:511];
  reg [63:0] GEN_9;
  wire [63:0] T_889_0_T_915_data;
  wire [8:0] T_889_0_T_915_addr;
  wire  T_889_0_T_915_en;
  reg [8:0] GEN_11;
  reg [31:0] GEN_12;
  reg  GEN_13;
  reg [31:0] GEN_14;
  wire [63:0] T_889_0_T_906_data;
  wire [8:0] T_889_0_T_906_addr;
  wire  T_889_0_T_906_mask;
  wire  T_889_0_T_906_en;
  wire  T_892;
  wire  T_894;
  wire [63:0] T_901_0;
  wire  GEN_18;
  wire [8:0] T_912;
  wire [63:0] T_923_0;
  wire  T_925;
  wire [63:0] T_933_0;
  reg [11:0] T_935;
  reg [31:0] GEN_15;
  wire [11:0] GEN_20;
  reg [63:0] T_944_0 [0:511];
  reg [63:0] GEN_16;
  wire [63:0] T_944_0_T_970_data;
  wire [8:0] T_944_0_T_970_addr;
  wire  T_944_0_T_970_en;
  reg [8:0] GEN_17;
  reg [31:0] GEN_19;
  reg  GEN_21;
  reg [31:0] GEN_22;
  wire [63:0] T_944_0_T_961_data;
  wire [8:0] T_944_0_T_961_addr;
  wire  T_944_0_T_961_mask;
  wire  T_944_0_T_961_en;
  wire  T_947;
  wire  T_949;
  wire [63:0] T_956_0;
  wire  GEN_28;
  wire [8:0] T_967;
  wire [63:0] T_978_0;
  wire  T_980;
  wire [63:0] T_988_0;
  reg [11:0] T_990;
  reg [31:0] GEN_23;
  wire [11:0] GEN_30;
  reg [63:0] T_999_0 [0:511];
  reg [63:0] GEN_24;
  wire [63:0] T_999_0_T_1025_data;
  wire [8:0] T_999_0_T_1025_addr;
  wire  T_999_0_T_1025_en;
  reg [8:0] GEN_25;
  reg [31:0] GEN_26;
  reg  GEN_27;
  reg [31:0] GEN_29;
  wire [63:0] T_999_0_T_1016_data;
  wire [8:0] T_999_0_T_1016_addr;
  wire  T_999_0_T_1016_mask;
  wire  T_999_0_T_1016_en;
  wire  T_1002;
  wire  T_1004;
  wire [63:0] T_1011_0;
  wire  GEN_38;
  wire [8:0] T_1022;
  wire [63:0] T_1033_0;
  assign io_read_ready = 1'h1;
  assign io_write_ready = 1'h1;
  assign io_resp_0 = T_868_0;
  assign io_resp_1 = T_923_0;
  assign io_resp_2 = T_978_0;
  assign io_resp_3 = T_1033_0;
  assign waddr = io_write_bits_addr[11:3];
  assign raddr = io_read_bits_addr[11:3];
  assign T_815 = io_write_bits_way_en[0];
  assign T_823_0 = T_834_0_T_860_data;
  assign GEN_0 = io_read_valid ? io_read_bits_addr : T_825;
  assign T_834_0_T_860_addr = T_857;
  assign T_834_0_T_860_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_834_0_T_860_data = T_834_0[GEN_3];
  `else
  assign T_834_0_T_860_data = GEN_3 >= 10'h200 ? $random : T_834_0[GEN_3];
  `endif
  assign T_834_0_T_851_data = T_846_0;
  assign T_834_0_T_851_addr = waddr;
  assign T_834_0_T_851_mask = GEN_8;
  assign T_834_0_T_851_en = T_839;
  assign T_837 = T_815 & io_write_valid;
  assign T_839 = T_837 & io_write_bits_wmask;
  assign T_846_0 = io_write_bits_data;
  assign GEN_8 = T_839 ? T_815 : 1'h0;
  assign T_857 = raddr;
  assign T_868_0 = T_823_0;
  assign T_870 = io_write_bits_way_en[1];
  assign T_878_0 = T_889_0_T_915_data;
  assign GEN_10 = io_read_valid ? io_read_bits_addr : T_880;
  assign T_889_0_T_915_addr = T_912;
  assign T_889_0_T_915_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_889_0_T_915_data = T_889_0[GEN_11];
  `else
  assign T_889_0_T_915_data = GEN_11 >= 10'h200 ? $random : T_889_0[GEN_11];
  `endif
  assign T_889_0_T_906_data = T_901_0;
  assign T_889_0_T_906_addr = waddr;
  assign T_889_0_T_906_mask = GEN_18;
  assign T_889_0_T_906_en = T_894;
  assign T_892 = T_870 & io_write_valid;
  assign T_894 = T_892 & io_write_bits_wmask;
  assign T_901_0 = io_write_bits_data;
  assign GEN_18 = T_894 ? T_870 : 1'h0;
  assign T_912 = raddr;
  assign T_923_0 = T_878_0;
  assign T_925 = io_write_bits_way_en[2];
  assign T_933_0 = T_944_0_T_970_data;
  assign GEN_20 = io_read_valid ? io_read_bits_addr : T_935;
  assign T_944_0_T_970_addr = T_967;
  assign T_944_0_T_970_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_944_0_T_970_data = T_944_0[GEN_17];
  `else
  assign T_944_0_T_970_data = GEN_17 >= 10'h200 ? $random : T_944_0[GEN_17];
  `endif
  assign T_944_0_T_961_data = T_956_0;
  assign T_944_0_T_961_addr = waddr;
  assign T_944_0_T_961_mask = GEN_28;
  assign T_944_0_T_961_en = T_949;
  assign T_947 = T_925 & io_write_valid;
  assign T_949 = T_947 & io_write_bits_wmask;
  assign T_956_0 = io_write_bits_data;
  assign GEN_28 = T_949 ? T_925 : 1'h0;
  assign T_967 = raddr;
  assign T_978_0 = T_933_0;
  assign T_980 = io_write_bits_way_en[3];
  assign T_988_0 = T_999_0_T_1025_data;
  assign GEN_30 = io_read_valid ? io_read_bits_addr : T_990;
  assign T_999_0_T_1025_addr = T_1022;
  assign T_999_0_T_1025_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_999_0_T_1025_data = T_999_0[GEN_25];
  `else
  assign T_999_0_T_1025_data = GEN_25 >= 10'h200 ? $random : T_999_0[GEN_25];
  `endif
  assign T_999_0_T_1016_data = T_1011_0;
  assign T_999_0_T_1016_addr = waddr;
  assign T_999_0_T_1016_mask = GEN_38;
  assign T_999_0_T_1016_en = T_1004;
  assign T_1002 = T_980 & io_write_valid;
  assign T_1004 = T_1002 & io_write_bits_wmask;
  assign T_1011_0 = io_write_bits_data;
  assign GEN_38 = T_1004 ? T_980 : 1'h0;
  assign T_1022 = raddr;
  assign T_1033_0 = T_988_0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_1 = {1{$random}};
  T_825 = GEN_1[11:0];
  GEN_2 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_834_0[initvar] = GEN_2[63:0];
  GEN_4 = {1{$random}};
  GEN_3 = GEN_4[8:0];
  GEN_6 = {1{$random}};
  GEN_5 = GEN_6[0:0];
  GEN_7 = {1{$random}};
  T_880 = GEN_7[11:0];
  GEN_9 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_889_0[initvar] = GEN_9[63:0];
  GEN_12 = {1{$random}};
  GEN_11 = GEN_12[8:0];
  GEN_14 = {1{$random}};
  GEN_13 = GEN_14[0:0];
  GEN_15 = {1{$random}};
  T_935 = GEN_15[11:0];
  GEN_16 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_944_0[initvar] = GEN_16[63:0];
  GEN_19 = {1{$random}};
  GEN_17 = GEN_19[8:0];
  GEN_22 = {1{$random}};
  GEN_21 = GEN_22[0:0];
  GEN_23 = {1{$random}};
  T_990 = GEN_23[11:0];
  GEN_24 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_999_0[initvar] = GEN_24[63:0];
  GEN_26 = {1{$random}};
  GEN_25 = GEN_26[8:0];
  GEN_29 = {1{$random}};
  GEN_27 = GEN_29[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(io_read_valid) begin
        T_825 <= io_read_bits_addr;
      end
    end
    GEN_3 <= T_834_0_T_860_addr;
    GEN_5 <= T_834_0_T_860_en;
    if(T_834_0_T_851_en & T_834_0_T_851_mask) begin
      T_834_0[T_834_0_T_851_addr] <= T_834_0_T_851_data;
    end
    if(1'h0) begin
    end else begin
      if(io_read_valid) begin
        T_880 <= io_read_bits_addr;
      end
    end
    GEN_11 <= T_889_0_T_915_addr;
    GEN_13 <= T_889_0_T_915_en;
    if(T_889_0_T_906_en & T_889_0_T_906_mask) begin
      T_889_0[T_889_0_T_906_addr] <= T_889_0_T_906_data;
    end
    if(1'h0) begin
    end else begin
      if(io_read_valid) begin
        T_935 <= io_read_bits_addr;
      end
    end
    GEN_17 <= T_944_0_T_970_addr;
    GEN_21 <= T_944_0_T_970_en;
    if(T_944_0_T_961_en & T_944_0_T_961_mask) begin
      T_944_0[T_944_0_T_961_addr] <= T_944_0_T_961_data;
    end
    if(1'h0) begin
    end else begin
      if(io_read_valid) begin
        T_990 <= io_read_bits_addr;
      end
    end
    GEN_25 <= T_999_0_T_1025_addr;
    GEN_27 <= T_999_0_T_1025_en;
    if(T_999_0_T_1016_en & T_999_0_T_1016_mask) begin
      T_999_0[T_999_0_T_1016_addr] <= T_999_0_T_1016_data;
    end
  end
endmodule
module Arbiter_10(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [3:0] io_in_0_bits_way_en,
  input  [11:0] io_in_0_bits_addr,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [3:0] io_in_1_bits_way_en,
  input  [11:0] io_in_1_bits_addr,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [3:0] io_in_2_bits_way_en,
  input  [11:0] io_in_2_bits_addr,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [3:0] io_in_3_bits_way_en,
  input  [11:0] io_in_3_bits_addr,
  input   io_out_ready,
  output  io_out_valid,
  output [3:0] io_out_bits_way_en,
  output [11:0] io_out_bits_addr,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [3:0] GEN_1;
  wire [11:0] GEN_2;
  wire [1:0] GEN_3;
  wire [3:0] GEN_4;
  wire [11:0] GEN_5;
  wire [1:0] GEN_6;
  wire [3:0] GEN_7;
  wire [11:0] GEN_8;
  wire  T_2205;
  wire  T_2206;
  wire  T_2208;
  wire  T_2210;
  wire  T_2212;
  wire  T_2214;
  wire  T_2215;
  wire  T_2216;
  wire  T_2218;
  wire  T_2219;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2214;
  assign io_in_2_ready = T_2215;
  assign io_in_3_ready = T_2216;
  assign io_out_valid = T_2219;
  assign io_out_bits_way_en = GEN_7;
  assign io_out_bits_addr = GEN_8;
  assign io_chosen = GEN_6;
  assign GEN_0 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_1 = io_in_2_valid ? io_in_2_bits_way_en : io_in_3_bits_way_en;
  assign GEN_2 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr;
  assign GEN_3 = io_in_1_valid ? {{1'd0}, 1'h1} : GEN_0;
  assign GEN_4 = io_in_1_valid ? io_in_1_bits_way_en : GEN_1;
  assign GEN_5 = io_in_1_valid ? io_in_1_bits_addr : GEN_2;
  assign GEN_6 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_3;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_way_en : GEN_4;
  assign GEN_8 = io_in_0_valid ? io_in_0_bits_addr : GEN_5;
  assign T_2205 = io_in_0_valid | io_in_1_valid;
  assign T_2206 = T_2205 | io_in_2_valid;
  assign T_2208 = io_in_0_valid == 1'h0;
  assign T_2210 = T_2205 == 1'h0;
  assign T_2212 = T_2206 == 1'h0;
  assign T_2214 = T_2208 & io_out_ready;
  assign T_2215 = T_2210 & io_out_ready;
  assign T_2216 = T_2212 & io_out_ready;
  assign T_2218 = T_2212 == 1'h0;
  assign T_2219 = T_2218 | io_in_3_valid;
endmodule
module Arbiter_11(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [3:0] io_in_0_bits_way_en,
  input  [11:0] io_in_0_bits_addr,
  input   io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [3:0] io_in_1_bits_way_en,
  input  [11:0] io_in_1_bits_addr,
  input   io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [3:0] io_out_bits_way_en,
  output [11:0] io_out_bits_addr,
  output  io_out_bits_wmask,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  GEN_0;
  wire [3:0] GEN_1;
  wire [11:0] GEN_2;
  wire  GEN_3;
  wire [63:0] GEN_4;
  wire  T_1664;
  wire  T_1666;
  wire  T_1668;
  wire  T_1669;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1666;
  assign io_out_valid = T_1669;
  assign io_out_bits_way_en = GEN_1;
  assign io_out_bits_addr = GEN_2;
  assign io_out_bits_wmask = GEN_3;
  assign io_out_bits_data = GEN_4;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_wmask : io_in_1_bits_wmask;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign T_1664 = io_in_0_valid == 1'h0;
  assign T_1666 = T_1664 & io_out_ready;
  assign T_1668 = T_1664 == 1'h0;
  assign T_1669 = T_1668 | io_in_1_valid;
endmodule
module AMOALU(
  input   clk,
  input   reset,
  input  [5:0] io_addr,
  input  [4:0] io_cmd,
  input  [2:0] io_typ,
  input  [63:0] io_lhs,
  input  [63:0] io_rhs,
  output [63:0] io_out
);
  wire [1:0] T_6;
  wire  T_8;
  wire [31:0] T_9;
  wire [63:0] T_10;
  wire [63:0] rhs;
  wire  T_11;
  wire  T_12;
  wire  sgned;
  wire  T_14;
  wire  max;
  wire  T_16;
  wire  min;
  wire  T_17;
  wire  T_18;
  wire  T_19;
  wire  T_20;
  wire  T_21;
  wire  T_22;
  wire  word;
  wire  T_25;
  wire [31:0] GEN_0;
  wire [31:0] T_26;
  wire [63:0] GEN_1;
  wire [63:0] T_27;
  wire [63:0] T_28;
  wire [63:0] T_29;
  wire [64:0] T_30;
  wire [63:0] adder_out;
  wire  T_33;
  wire  T_34;
  wire  T_35;
  wire  T_36;
  wire  T_37;
  wire  T_42;
  wire  T_43;
  wire  T_44;
  wire [31:0] T_45;
  wire [31:0] T_46;
  wire  T_47;
  wire [31:0] T_48;
  wire [31:0] T_49;
  wire  T_50;
  wire  T_53;
  wire  T_55;
  wire  T_56;
  wire  T_57;
  wire  T_58;
  wire  T_59;
  wire  T_60;
  wire  less;
  wire  T_61;
  wire  T_62;
  wire [63:0] T_63;
  wire  T_64;
  wire [63:0] T_65;
  wire  T_66;
  wire [63:0] T_67;
  wire  T_68;
  wire [1:0] GEN_2;
  wire  T_70;
  wire [7:0] T_71;
  wire [15:0] T_72;
  wire [31:0] T_73;
  wire [63:0] T_74;
  wire [1:0] GEN_3;
  wire  T_76;
  wire [15:0] T_77;
  wire [31:0] T_78;
  wire [63:0] T_79;
  wire [63:0] T_85;
  wire [63:0] T_86;
  wire [63:0] T_87;
  wire [63:0] T_88;
  wire [63:0] T_89;
  wire [63:0] T_90;
  wire [63:0] out;
  wire  T_92;
  wire  T_96;
  wire  T_100;
  wire  T_103;
  wire [1:0] T_104;
  wire  T_105;
  wire [1:0] T_107;
  wire  T_109;
  wire [1:0] T_112;
  wire [1:0] T_113;
  wire [1:0] T_116;
  wire [3:0] T_117;
  wire [3:0] T_120;
  wire  T_122;
  wire [3:0] T_125;
  wire [3:0] T_126;
  wire [3:0] T_129;
  wire [7:0] T_130;
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire  T_134;
  wire  T_135;
  wire  T_136;
  wire  T_137;
  wire  T_138;
  wire [7:0] GEN_5;
  wire [8:0] T_140;
  wire [7:0] T_141;
  wire [7:0] GEN_6;
  wire [8:0] T_143;
  wire [7:0] T_144;
  wire [7:0] GEN_7;
  wire [8:0] T_146;
  wire [7:0] T_147;
  wire [7:0] GEN_8;
  wire [8:0] T_149;
  wire [7:0] T_150;
  wire [7:0] GEN_9;
  wire [8:0] T_152;
  wire [7:0] T_153;
  wire [7:0] GEN_10;
  wire [8:0] T_155;
  wire [7:0] T_156;
  wire [7:0] GEN_11;
  wire [8:0] T_158;
  wire [7:0] T_159;
  wire [7:0] GEN_12;
  wire [8:0] T_161;
  wire [7:0] T_162;
  wire [7:0] T_168_0;
  wire [7:0] T_168_1;
  wire [7:0] T_168_2;
  wire [7:0] T_168_3;
  wire [7:0] T_168_4;
  wire [7:0] T_168_5;
  wire [7:0] T_168_6;
  wire [7:0] T_168_7;
  wire [15:0] T_170;
  wire [15:0] T_171;
  wire [31:0] T_172;
  wire [15:0] T_173;
  wire [15:0] T_174;
  wire [31:0] T_175;
  wire [63:0] wmask;
  wire [63:0] T_176;
  wire [63:0] T_177;
  wire [63:0] T_178;
  wire [63:0] T_179;
  assign io_out = T_179;
  assign T_6 = io_typ[1:0];
  assign T_8 = T_6 == 2'h2;
  assign T_9 = io_rhs[31:0];
  assign T_10 = {T_9,T_9};
  assign rhs = T_8 ? T_10 : io_rhs;
  assign T_11 = io_cmd == 5'hc;
  assign T_12 = io_cmd == 5'hd;
  assign sgned = T_11 | T_12;
  assign T_14 = io_cmd == 5'hf;
  assign max = T_12 | T_14;
  assign T_16 = io_cmd == 5'he;
  assign min = T_11 | T_16;
  assign T_17 = io_typ == 3'h2;
  assign T_18 = io_typ == 3'h6;
  assign T_19 = T_17 | T_18;
  assign T_20 = io_typ == 3'h0;
  assign T_21 = T_19 | T_20;
  assign T_22 = io_typ == 3'h4;
  assign word = T_21 | T_22;
  assign T_25 = io_addr[2];
  assign GEN_0 = {{31'd0}, T_25};
  assign T_26 = GEN_0 << 31;
  assign GEN_1 = {{32'd0}, T_26};
  assign T_27 = 64'hffffffffffffffff ^ GEN_1;
  assign T_28 = io_lhs & T_27;
  assign T_29 = rhs & T_27;
  assign T_30 = T_28 + T_29;
  assign adder_out = T_30[63:0];
  assign T_33 = T_25 == 1'h0;
  assign T_34 = word & T_33;
  assign T_35 = io_lhs[31];
  assign T_36 = io_lhs[63];
  assign T_37 = T_34 ? T_35 : T_36;
  assign T_42 = rhs[31];
  assign T_43 = rhs[63];
  assign T_44 = T_34 ? T_42 : T_43;
  assign T_45 = io_lhs[31:0];
  assign T_46 = rhs[31:0];
  assign T_47 = T_45 < T_46;
  assign T_48 = io_lhs[63:32];
  assign T_49 = rhs[63:32];
  assign T_50 = T_48 < T_49;
  assign T_53 = T_48 == T_49;
  assign T_55 = T_25 ? T_50 : T_47;
  assign T_56 = T_53 & T_47;
  assign T_57 = T_50 | T_56;
  assign T_58 = word ? T_55 : T_57;
  assign T_59 = T_37 == T_44;
  assign T_60 = sgned ? T_37 : T_44;
  assign less = T_59 ? T_58 : T_60;
  assign T_61 = io_cmd == 5'h8;
  assign T_62 = io_cmd == 5'hb;
  assign T_63 = io_lhs & rhs;
  assign T_64 = io_cmd == 5'ha;
  assign T_65 = io_lhs | rhs;
  assign T_66 = io_cmd == 5'h9;
  assign T_67 = io_lhs ^ rhs;
  assign T_68 = less ? min : max;
  assign GEN_2 = {{1'd0}, 1'h0};
  assign T_70 = T_6 == GEN_2;
  assign T_71 = io_rhs[7:0];
  assign T_72 = {T_71,T_71};
  assign T_73 = {T_72,T_72};
  assign T_74 = {T_73,T_73};
  assign GEN_3 = {{1'd0}, 1'h1};
  assign T_76 = T_6 == GEN_3;
  assign T_77 = io_rhs[15:0];
  assign T_78 = {T_77,T_77};
  assign T_79 = {T_78,T_78};
  assign T_85 = T_76 ? T_79 : rhs;
  assign T_86 = T_70 ? T_74 : T_85;
  assign T_87 = T_68 ? io_lhs : T_86;
  assign T_88 = T_66 ? T_67 : T_87;
  assign T_89 = T_64 ? T_65 : T_88;
  assign T_90 = T_62 ? T_63 : T_89;
  assign out = T_61 ? adder_out : T_90;
  assign T_92 = io_addr[0];
  assign T_96 = T_6 >= GEN_3;
  assign T_100 = T_92 | T_96;
  assign T_103 = T_92 ? 1'h0 : 1'h1;
  assign T_104 = {T_100,T_103};
  assign T_105 = io_addr[1];
  assign T_107 = T_105 ? T_104 : {{1'd0}, 1'h0};
  assign T_109 = T_6 >= 2'h2;
  assign T_112 = T_109 ? 2'h3 : {{1'd0}, 1'h0};
  assign T_113 = T_107 | T_112;
  assign T_116 = T_105 ? {{1'd0}, 1'h0} : T_104;
  assign T_117 = {T_113,T_116};
  assign T_120 = T_25 ? T_117 : {{3'd0}, 1'h0};
  assign T_122 = T_6 >= 2'h3;
  assign T_125 = T_122 ? 4'hf : {{3'd0}, 1'h0};
  assign T_126 = T_120 | T_125;
  assign T_129 = T_25 ? {{3'd0}, 1'h0} : T_117;
  assign T_130 = {T_126,T_129};
  assign T_131 = T_130[0];
  assign T_132 = T_130[1];
  assign T_133 = T_130[2];
  assign T_134 = T_130[3];
  assign T_135 = T_130[4];
  assign T_136 = T_130[5];
  assign T_137 = T_130[6];
  assign T_138 = T_130[7];
  assign GEN_5 = {{7'd0}, T_131};
  assign T_140 = 8'h0 - GEN_5;
  assign T_141 = T_140[7:0];
  assign GEN_6 = {{7'd0}, T_132};
  assign T_143 = 8'h0 - GEN_6;
  assign T_144 = T_143[7:0];
  assign GEN_7 = {{7'd0}, T_133};
  assign T_146 = 8'h0 - GEN_7;
  assign T_147 = T_146[7:0];
  assign GEN_8 = {{7'd0}, T_134};
  assign T_149 = 8'h0 - GEN_8;
  assign T_150 = T_149[7:0];
  assign GEN_9 = {{7'd0}, T_135};
  assign T_152 = 8'h0 - GEN_9;
  assign T_153 = T_152[7:0];
  assign GEN_10 = {{7'd0}, T_136};
  assign T_155 = 8'h0 - GEN_10;
  assign T_156 = T_155[7:0];
  assign GEN_11 = {{7'd0}, T_137};
  assign T_158 = 8'h0 - GEN_11;
  assign T_159 = T_158[7:0];
  assign GEN_12 = {{7'd0}, T_138};
  assign T_161 = 8'h0 - GEN_12;
  assign T_162 = T_161[7:0];
  assign T_168_0 = T_141;
  assign T_168_1 = T_144;
  assign T_168_2 = T_147;
  assign T_168_3 = T_150;
  assign T_168_4 = T_153;
  assign T_168_5 = T_156;
  assign T_168_6 = T_159;
  assign T_168_7 = T_162;
  assign T_170 = {T_168_1,T_168_0};
  assign T_171 = {T_168_3,T_168_2};
  assign T_172 = {T_171,T_170};
  assign T_173 = {T_168_5,T_168_4};
  assign T_174 = {T_168_7,T_168_6};
  assign T_175 = {T_174,T_173};
  assign wmask = {T_175,T_172};
  assign T_176 = wmask & out;
  assign T_177 = ~ wmask;
  assign T_178 = T_177 & io_lhs;
  assign T_179 = T_176 | T_178;
endmodule
module LockingArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_7;
  wire [2:0] GEN_1;
  wire [2:0] GEN_8;
  wire [25:0] GEN_2;
  wire [25:0] GEN_9;
  wire [1:0] GEN_3;
  wire [1:0] GEN_10;
  wire  GEN_4;
  wire  GEN_11;
  wire [2:0] GEN_5;
  wire [2:0] GEN_12;
  wire [63:0] GEN_6;
  wire [63:0] GEN_13;
  reg [2:0] T_818;
  reg [31:0] GEN_20;
  reg  T_820;
  reg [31:0] GEN_21;
  wire [2:0] GEN_18;
  wire  T_822;
  wire [2:0] T_829_0;
  wire [2:0] T_829_1;
  wire [2:0] T_829_2;
  wire  T_831;
  wire  T_832;
  wire  T_833;
  wire  T_836;
  wire  T_837;
  wire  T_839;
  wire  T_840;
  wire [2:0] GEN_19;
  wire [3:0] T_844;
  wire [2:0] T_845;
  wire  GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  wire  T_848;
  wire  T_850;
  wire  T_851;
  wire  T_852;
  wire  T_855;
  wire  T_856;
  wire  GEN_17;
  assign io_in_0_ready = T_852;
  assign io_in_1_ready = T_856;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_addr_block = GEN_2;
  assign io_out_bits_client_xact_id = GEN_3;
  assign io_out_bits_voluntary = GEN_4;
  assign io_out_bits_r_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_16;
  assign choice = GEN_17;
  assign GEN_0 = GEN_7;
  assign GEN_7 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_2 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_3 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_4 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign GEN_5 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign GEN_6 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_18 = {{2'd0}, 1'h0};
  assign T_822 = T_818 != GEN_18;
  assign T_829_0 = 3'h0;
  assign T_829_1 = 3'h1;
  assign T_829_2 = 3'h2;
  assign T_831 = T_829_0 == io_out_bits_r_type;
  assign T_832 = T_829_1 == io_out_bits_r_type;
  assign T_833 = T_829_2 == io_out_bits_r_type;
  assign T_836 = T_831 | T_832;
  assign T_837 = T_836 | T_833;
  assign T_839 = io_out_ready & io_out_valid;
  assign T_840 = T_839 & T_837;
  assign GEN_19 = {{2'd0}, 1'h1};
  assign T_844 = T_818 + GEN_19;
  assign T_845 = T_844[2:0];
  assign GEN_14 = T_840 ? io_chosen : T_820;
  assign GEN_15 = T_840 ? T_845 : T_818;
  assign GEN_16 = T_822 ? T_820 : choice;
  assign T_848 = io_in_0_valid == 1'h0;
  assign T_850 = T_820 == 1'h0;
  assign T_851 = T_822 ? T_850 : 1'h1;
  assign T_852 = T_851 & io_out_ready;
  assign T_855 = T_822 ? T_820 : T_848;
  assign T_856 = T_855 & io_out_ready;
  assign GEN_17 = io_in_0_valid ? 1'h0 : 1'h1;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_20 = {1{$random}};
  T_818 = GEN_20[2:0];
  GEN_21 = {1{$random}};
  T_820 = GEN_21[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_818 <= 3'h0;
    end else begin
      if(T_840) begin
        T_818 <= T_845;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_840) begin
        T_820 <= io_chosen;
      end
    end
  end
endmodule
module FlowThroughSerializer_1(
  input   clk,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input  [2:0] io_in_bits_addr_beat,
  input  [1:0] io_in_bits_client_xact_id,
  input  [2:0] io_in_bits_manager_xact_id,
  input   io_in_bits_is_builtin_type,
  input  [3:0] io_in_bits_g_type,
  input  [63:0] io_in_bits_data,
  input   io_in_bits_manager_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_manager_id,
  output  io_cnt,
  output  io_done
);
  assign io_in_ready = io_out_ready;
  assign io_out_valid = io_in_valid;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_data = io_in_bits_data;
  assign io_out_bits_manager_id = io_in_bits_manager_id;
  assign io_cnt = 1'h0;
  assign io_done = 1'h1;
endmodule
module HellaCache(
  input   clk,
  input   reset,
  output  io_cpu_req_ready,
  input   io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_addr,
  input  [8:0] io_cpu_req_bits_tag,
  input  [4:0] io_cpu_req_bits_cmd,
  input  [2:0] io_cpu_req_bits_typ,
  input   io_cpu_req_bits_phys,
  input  [63:0] io_cpu_req_bits_data,
  input   io_cpu_s1_kill,
  input  [63:0] io_cpu_s1_data,
  output  io_cpu_s2_nack,
  output  io_cpu_resp_valid,
  output [39:0] io_cpu_resp_bits_addr,
  output [8:0] io_cpu_resp_bits_tag,
  output [4:0] io_cpu_resp_bits_cmd,
  output [2:0] io_cpu_resp_bits_typ,
  output [63:0] io_cpu_resp_bits_data,
  output  io_cpu_resp_bits_replay,
  output  io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output [63:0] io_cpu_resp_bits_store_data,
  output  io_cpu_replay_next,
  output  io_cpu_xcpt_ma_ld,
  output  io_cpu_xcpt_ma_st,
  output  io_cpu_xcpt_pf_ld,
  output  io_cpu_xcpt_pf_st,
  input   io_cpu_invalidate_lr,
  output  io_cpu_ordered,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_addr,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [19:0] io_ptw_resp_bits_pte_ppn,
  input  [2:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_r,
  input  [3:0] io_ptw_resp_bits_pte_typ,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [4:0] io_ptw_status_zero1,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_probe_ready,
  input   io_mem_probe_valid,
  input  [25:0] io_mem_probe_bits_addr_block,
  input  [1:0] io_mem_probe_bits_p_type,
  input   io_mem_release_ready,
  output  io_mem_release_valid,
  output [2:0] io_mem_release_bits_addr_beat,
  output [25:0] io_mem_release_bits_addr_block,
  output [1:0] io_mem_release_bits_client_xact_id,
  output  io_mem_release_bits_voluntary,
  output [2:0] io_mem_release_bits_r_type,
  output [63:0] io_mem_release_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id
);
  wire  wb_clk;
  wire  wb_reset;
  wire  wb_io_req_ready;
  wire  wb_io_req_valid;
  wire [2:0] wb_io_req_bits_addr_beat;
  wire [25:0] wb_io_req_bits_addr_block;
  wire [1:0] wb_io_req_bits_client_xact_id;
  wire  wb_io_req_bits_voluntary;
  wire [2:0] wb_io_req_bits_r_type;
  wire [63:0] wb_io_req_bits_data;
  wire [3:0] wb_io_req_bits_way_en;
  wire  wb_io_meta_read_ready;
  wire  wb_io_meta_read_valid;
  wire [5:0] wb_io_meta_read_bits_idx;
  wire [3:0] wb_io_meta_read_bits_way_en;
  wire [19:0] wb_io_meta_read_bits_tag;
  wire  wb_io_data_req_ready;
  wire  wb_io_data_req_valid;
  wire [3:0] wb_io_data_req_bits_way_en;
  wire [11:0] wb_io_data_req_bits_addr;
  wire [63:0] wb_io_data_resp;
  wire  wb_io_release_ready;
  wire  wb_io_release_valid;
  wire [2:0] wb_io_release_bits_addr_beat;
  wire [25:0] wb_io_release_bits_addr_block;
  wire [1:0] wb_io_release_bits_client_xact_id;
  wire  wb_io_release_bits_voluntary;
  wire [2:0] wb_io_release_bits_r_type;
  wire [63:0] wb_io_release_bits_data;
  wire  prober_clk;
  wire  prober_reset;
  wire  prober_io_req_ready;
  wire  prober_io_req_valid;
  wire [25:0] prober_io_req_bits_addr_block;
  wire [1:0] prober_io_req_bits_p_type;
  wire [1:0] prober_io_req_bits_client_xact_id;
  wire  prober_io_rep_ready;
  wire  prober_io_rep_valid;
  wire [2:0] prober_io_rep_bits_addr_beat;
  wire [25:0] prober_io_rep_bits_addr_block;
  wire [1:0] prober_io_rep_bits_client_xact_id;
  wire  prober_io_rep_bits_voluntary;
  wire [2:0] prober_io_rep_bits_r_type;
  wire [63:0] prober_io_rep_bits_data;
  wire  prober_io_meta_read_ready;
  wire  prober_io_meta_read_valid;
  wire [5:0] prober_io_meta_read_bits_idx;
  wire [3:0] prober_io_meta_read_bits_way_en;
  wire [19:0] prober_io_meta_read_bits_tag;
  wire  prober_io_meta_write_ready;
  wire  prober_io_meta_write_valid;
  wire [5:0] prober_io_meta_write_bits_idx;
  wire [3:0] prober_io_meta_write_bits_way_en;
  wire [19:0] prober_io_meta_write_bits_data_tag;
  wire [1:0] prober_io_meta_write_bits_data_coh_state;
  wire  prober_io_wb_req_ready;
  wire  prober_io_wb_req_valid;
  wire [2:0] prober_io_wb_req_bits_addr_beat;
  wire [25:0] prober_io_wb_req_bits_addr_block;
  wire [1:0] prober_io_wb_req_bits_client_xact_id;
  wire  prober_io_wb_req_bits_voluntary;
  wire [2:0] prober_io_wb_req_bits_r_type;
  wire [63:0] prober_io_wb_req_bits_data;
  wire [3:0] prober_io_wb_req_bits_way_en;
  wire [3:0] prober_io_way_en;
  wire  prober_io_mshr_rdy;
  wire [1:0] prober_io_block_state_state;
  wire  mshrs_clk;
  wire  mshrs_reset;
  wire  mshrs_io_req_ready;
  wire  mshrs_io_req_valid;
  wire [39:0] mshrs_io_req_bits_addr;
  wire [8:0] mshrs_io_req_bits_tag;
  wire [4:0] mshrs_io_req_bits_cmd;
  wire [2:0] mshrs_io_req_bits_typ;
  wire  mshrs_io_req_bits_phys;
  wire [63:0] mshrs_io_req_bits_data;
  wire  mshrs_io_req_bits_tag_match;
  wire [19:0] mshrs_io_req_bits_old_meta_tag;
  wire [1:0] mshrs_io_req_bits_old_meta_coh_state;
  wire [3:0] mshrs_io_req_bits_way_en;
  wire  mshrs_io_resp_ready;
  wire  mshrs_io_resp_valid;
  wire [39:0] mshrs_io_resp_bits_addr;
  wire [8:0] mshrs_io_resp_bits_tag;
  wire [4:0] mshrs_io_resp_bits_cmd;
  wire [2:0] mshrs_io_resp_bits_typ;
  wire [63:0] mshrs_io_resp_bits_data;
  wire  mshrs_io_resp_bits_replay;
  wire  mshrs_io_resp_bits_has_data;
  wire [63:0] mshrs_io_resp_bits_data_word_bypass;
  wire [63:0] mshrs_io_resp_bits_store_data;
  wire  mshrs_io_secondary_miss;
  wire  mshrs_io_mem_req_ready;
  wire  mshrs_io_mem_req_valid;
  wire [25:0] mshrs_io_mem_req_bits_addr_block;
  wire [1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire [2:0] mshrs_io_mem_req_bits_addr_beat;
  wire  mshrs_io_mem_req_bits_is_builtin_type;
  wire [2:0] mshrs_io_mem_req_bits_a_type;
  wire [11:0] mshrs_io_mem_req_bits_union;
  wire [63:0] mshrs_io_mem_req_bits_data;
  wire [3:0] mshrs_io_refill_way_en;
  wire [11:0] mshrs_io_refill_addr;
  wire  mshrs_io_meta_read_ready;
  wire  mshrs_io_meta_read_valid;
  wire [5:0] mshrs_io_meta_read_bits_idx;
  wire [3:0] mshrs_io_meta_read_bits_way_en;
  wire [19:0] mshrs_io_meta_read_bits_tag;
  wire  mshrs_io_meta_write_ready;
  wire  mshrs_io_meta_write_valid;
  wire [5:0] mshrs_io_meta_write_bits_idx;
  wire [3:0] mshrs_io_meta_write_bits_way_en;
  wire [19:0] mshrs_io_meta_write_bits_data_tag;
  wire [1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire  mshrs_io_replay_ready;
  wire  mshrs_io_replay_valid;
  wire [39:0] mshrs_io_replay_bits_addr;
  wire [8:0] mshrs_io_replay_bits_tag;
  wire [4:0] mshrs_io_replay_bits_cmd;
  wire [2:0] mshrs_io_replay_bits_typ;
  wire  mshrs_io_replay_bits_phys;
  wire [63:0] mshrs_io_replay_bits_data;
  wire  mshrs_io_mem_grant_valid;
  wire [2:0] mshrs_io_mem_grant_bits_addr_beat;
  wire [1:0] mshrs_io_mem_grant_bits_client_xact_id;
  wire [2:0] mshrs_io_mem_grant_bits_manager_xact_id;
  wire  mshrs_io_mem_grant_bits_is_builtin_type;
  wire [3:0] mshrs_io_mem_grant_bits_g_type;
  wire [63:0] mshrs_io_mem_grant_bits_data;
  wire  mshrs_io_mem_grant_bits_manager_id;
  wire  mshrs_io_mem_finish_ready;
  wire  mshrs_io_mem_finish_valid;
  wire [2:0] mshrs_io_mem_finish_bits_manager_xact_id;
  wire  mshrs_io_mem_finish_bits_manager_id;
  wire  mshrs_io_wb_req_ready;
  wire  mshrs_io_wb_req_valid;
  wire [2:0] mshrs_io_wb_req_bits_addr_beat;
  wire [25:0] mshrs_io_wb_req_bits_addr_block;
  wire [1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire  mshrs_io_wb_req_bits_voluntary;
  wire [2:0] mshrs_io_wb_req_bits_r_type;
  wire [63:0] mshrs_io_wb_req_bits_data;
  wire [3:0] mshrs_io_wb_req_bits_way_en;
  wire  mshrs_io_probe_rdy;
  wire  mshrs_io_fence_rdy;
  wire  mshrs_io_replay_next;
  wire  T_2081;
  reg  s1_valid;
  reg [31:0] GEN_94;
  reg [39:0] s1_req_addr;
  reg [63:0] GEN_104;
  reg [8:0] s1_req_tag;
  reg [31:0] GEN_105;
  reg [4:0] s1_req_cmd;
  reg [31:0] GEN_109;
  reg [2:0] s1_req_typ;
  reg [31:0] GEN_114;
  reg  s1_req_phys;
  reg [31:0] GEN_115;
  reg [63:0] s1_req_data;
  reg [63:0] GEN_116;
  wire  T_2159;
  wire  s1_valid_masked;
  reg  s1_replay;
  reg [31:0] GEN_117;
  reg  s1_clk_en;
  reg [31:0] GEN_118;
  reg  s2_valid;
  reg [31:0] GEN_119;
  reg [39:0] s2_req_addr;
  reg [63:0] GEN_120;
  reg [8:0] s2_req_tag;
  reg [31:0] GEN_121;
  reg [4:0] s2_req_cmd;
  reg [31:0] GEN_122;
  reg [2:0] s2_req_typ;
  reg [31:0] GEN_123;
  reg  s2_req_phys;
  reg [31:0] GEN_124;
  reg [63:0] s2_req_data;
  reg [63:0] GEN_125;
  reg  T_2239;
  reg [31:0] GEN_126;
  wire  T_2240;
  wire  s2_replay;
  wire  s2_recycle;
  wire  s2_valid_masked;
  reg  s3_valid;
  reg [31:0] GEN_127;
  reg [39:0] s3_req_addr;
  reg [63:0] GEN_128;
  reg [8:0] s3_req_tag;
  reg [31:0] GEN_129;
  reg [4:0] s3_req_cmd;
  reg [31:0] GEN_130;
  reg [2:0] s3_req_typ;
  reg [31:0] GEN_131;
  reg  s3_req_phys;
  reg [31:0] GEN_132;
  reg [63:0] s3_req_data;
  reg [63:0] GEN_133;
  reg [3:0] s3_way;
  reg [31:0] GEN_134;
  reg  s1_recycled;
  reg [31:0] GEN_135;
  wire  GEN_0;
  wire  T_2321;
  wire  T_2322;
  wire  T_2323;
  wire  T_2324;
  wire  T_2325;
  wire  T_2326;
  wire  T_2327;
  wire  T_2328;
  wire  s1_read;
  wire  T_2329;
  wire  T_2331;
  wire  s1_write;
  wire  T_2335;
  wire  T_2336;
  wire  T_2337;
  wire  T_2338;
  wire  s1_readwrite;
  wire  dtlb_clk;
  wire  dtlb_reset;
  wire  dtlb_io_req_ready;
  wire  dtlb_io_req_valid;
  wire [27:0] dtlb_io_req_bits_vpn;
  wire  dtlb_io_req_bits_passthrough;
  wire  dtlb_io_req_bits_instruction;
  wire  dtlb_io_req_bits_store;
  wire  dtlb_io_resp_miss;
  wire [19:0] dtlb_io_resp_ppn;
  wire  dtlb_io_resp_xcpt_ld;
  wire  dtlb_io_resp_xcpt_st;
  wire  dtlb_io_resp_xcpt_if;
  wire [7:0] dtlb_io_resp_hit_idx;
  wire  dtlb_io_ptw_req_ready;
  wire  dtlb_io_ptw_req_valid;
  wire [26:0] dtlb_io_ptw_req_bits_addr;
  wire [1:0] dtlb_io_ptw_req_bits_prv;
  wire  dtlb_io_ptw_req_bits_store;
  wire  dtlb_io_ptw_req_bits_fetch;
  wire  dtlb_io_ptw_resp_valid;
  wire [19:0] dtlb_io_ptw_resp_bits_pte_ppn;
  wire [2:0] dtlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  dtlb_io_ptw_resp_bits_pte_d;
  wire  dtlb_io_ptw_resp_bits_pte_r;
  wire [3:0] dtlb_io_ptw_resp_bits_pte_typ;
  wire  dtlb_io_ptw_resp_bits_pte_v;
  wire [6:0] dtlb_io_ptw_ptbr_asid;
  wire [37:0] dtlb_io_ptw_ptbr_ppn;
  wire  dtlb_io_ptw_invalidate;
  wire  dtlb_io_ptw_status_debug;
  wire [1:0] dtlb_io_ptw_status_prv;
  wire  dtlb_io_ptw_status_sd;
  wire [30:0] dtlb_io_ptw_status_zero3;
  wire  dtlb_io_ptw_status_sd_rv32;
  wire [1:0] dtlb_io_ptw_status_zero2;
  wire [4:0] dtlb_io_ptw_status_vm;
  wire [4:0] dtlb_io_ptw_status_zero1;
  wire  dtlb_io_ptw_status_pum;
  wire  dtlb_io_ptw_status_mprv;
  wire [1:0] dtlb_io_ptw_status_xs;
  wire [1:0] dtlb_io_ptw_status_fs;
  wire [1:0] dtlb_io_ptw_status_mpp;
  wire [1:0] dtlb_io_ptw_status_hpp;
  wire  dtlb_io_ptw_status_spp;
  wire  dtlb_io_ptw_status_mpie;
  wire  dtlb_io_ptw_status_hpie;
  wire  dtlb_io_ptw_status_spie;
  wire  dtlb_io_ptw_status_upie;
  wire  dtlb_io_ptw_status_mie;
  wire  dtlb_io_ptw_status_hie;
  wire  dtlb_io_ptw_status_sie;
  wire  dtlb_io_ptw_status_uie;
  wire  T_2339;
  wire [27:0] T_2340;
  wire  T_2343;
  wire  T_2345;
  wire  T_2346;
  wire  GEN_1;
  wire [39:0] GEN_2;
  wire [8:0] GEN_3;
  wire [4:0] GEN_4;
  wire [2:0] GEN_5;
  wire  GEN_6;
  wire [63:0] GEN_7;
  wire [25:0] T_2348;
  wire [31:0] GEN_83;
  wire [31:0] T_2349;
  wire [39:0] GEN_8;
  wire  GEN_9;
  wire [25:0] T_2351;
  wire [31:0] GEN_84;
  wire [31:0] T_2352;
  wire [39:0] GEN_10;
  wire  GEN_11;
  wire [39:0] GEN_12;
  wire [8:0] GEN_13;
  wire [4:0] GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  wire [63:0] GEN_17;
  wire [39:0] GEN_18;
  wire [8:0] GEN_19;
  wire [4:0] GEN_20;
  wire [2:0] GEN_21;
  wire  GEN_22;
  wire [63:0] GEN_23;
  wire [11:0] T_2354;
  wire [31:0] s1_addr;
  wire [63:0] T_2355;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [2:0] GEN_26;
  wire  GEN_27;
  wire [39:0] GEN_28;
  wire [63:0] GEN_29;
  wire [8:0] GEN_30;
  wire [4:0] GEN_31;
  wire [1:0] T_2357;
  wire [3:0] GEN_85;
  wire [3:0] T_2359;
  wire [4:0] T_2361;
  wire [3:0] T_2362;
  wire [2:0] T_2363;
  wire [39:0] GEN_87;
  wire [39:0] T_2364;
  wire [39:0] GEN_88;
  wire  misaligned;
  wire  T_2366;
  wire  T_2367;
  wire  T_2368;
  wire  T_2369;
  wire  T_2370;
  wire  T_2371;
  wire  T_2372;
  reg  T_2373;
  reg [31:0] GEN_136;
  wire  T_2374;
  wire  T_2376;
  wire  T_2377;
  wire  T_2379;
  wire  meta_clk;
  wire  meta_reset;
  wire  meta_io_read_ready;
  wire  meta_io_read_valid;
  wire [5:0] meta_io_read_bits_idx;
  wire [3:0] meta_io_read_bits_way_en;
  wire  meta_io_write_ready;
  wire  meta_io_write_valid;
  wire [5:0] meta_io_write_bits_idx;
  wire [3:0] meta_io_write_bits_way_en;
  wire [19:0] meta_io_write_bits_data_tag;
  wire [1:0] meta_io_write_bits_data_coh_state;
  wire [19:0] meta_io_resp_0_tag;
  wire [1:0] meta_io_resp_0_coh_state;
  wire [19:0] meta_io_resp_1_tag;
  wire [1:0] meta_io_resp_1_coh_state;
  wire [19:0] meta_io_resp_2_tag;
  wire [1:0] meta_io_resp_2_coh_state;
  wire [19:0] meta_io_resp_3_tag;
  wire [1:0] meta_io_resp_3_coh_state;
  wire  metaReadArb_clk;
  wire  metaReadArb_reset;
  wire  metaReadArb_io_in_0_ready;
  wire  metaReadArb_io_in_0_valid;
  wire [5:0] metaReadArb_io_in_0_bits_idx;
  wire [3:0] metaReadArb_io_in_0_bits_way_en;
  wire  metaReadArb_io_in_1_ready;
  wire  metaReadArb_io_in_1_valid;
  wire [5:0] metaReadArb_io_in_1_bits_idx;
  wire [3:0] metaReadArb_io_in_1_bits_way_en;
  wire  metaReadArb_io_in_2_ready;
  wire  metaReadArb_io_in_2_valid;
  wire [5:0] metaReadArb_io_in_2_bits_idx;
  wire [3:0] metaReadArb_io_in_2_bits_way_en;
  wire  metaReadArb_io_in_3_ready;
  wire  metaReadArb_io_in_3_valid;
  wire [5:0] metaReadArb_io_in_3_bits_idx;
  wire [3:0] metaReadArb_io_in_3_bits_way_en;
  wire  metaReadArb_io_in_4_ready;
  wire  metaReadArb_io_in_4_valid;
  wire [5:0] metaReadArb_io_in_4_bits_idx;
  wire [3:0] metaReadArb_io_in_4_bits_way_en;
  wire  metaReadArb_io_out_ready;
  wire  metaReadArb_io_out_valid;
  wire [5:0] metaReadArb_io_out_bits_idx;
  wire [3:0] metaReadArb_io_out_bits_way_en;
  wire [2:0] metaReadArb_io_chosen;
  wire  metaWriteArb_clk;
  wire  metaWriteArb_reset;
  wire  metaWriteArb_io_in_0_ready;
  wire  metaWriteArb_io_in_0_valid;
  wire [5:0] metaWriteArb_io_in_0_bits_idx;
  wire [3:0] metaWriteArb_io_in_0_bits_way_en;
  wire [19:0] metaWriteArb_io_in_0_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_0_bits_data_coh_state;
  wire  metaWriteArb_io_in_1_ready;
  wire  metaWriteArb_io_in_1_valid;
  wire [5:0] metaWriteArb_io_in_1_bits_idx;
  wire [3:0] metaWriteArb_io_in_1_bits_way_en;
  wire [19:0] metaWriteArb_io_in_1_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_1_bits_data_coh_state;
  wire  metaWriteArb_io_out_ready;
  wire  metaWriteArb_io_out_valid;
  wire [5:0] metaWriteArb_io_out_bits_idx;
  wire [3:0] metaWriteArb_io_out_bits_way_en;
  wire [19:0] metaWriteArb_io_out_bits_data_tag;
  wire [1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire  metaWriteArb_io_chosen;
  wire  data_clk;
  wire  data_reset;
  wire  data_io_read_ready;
  wire  data_io_read_valid;
  wire [3:0] data_io_read_bits_way_en;
  wire [11:0] data_io_read_bits_addr;
  wire  data_io_write_ready;
  wire  data_io_write_valid;
  wire [3:0] data_io_write_bits_way_en;
  wire [11:0] data_io_write_bits_addr;
  wire  data_io_write_bits_wmask;
  wire [63:0] data_io_write_bits_data;
  wire [63:0] data_io_resp_0;
  wire [63:0] data_io_resp_1;
  wire [63:0] data_io_resp_2;
  wire [63:0] data_io_resp_3;
  wire  readArb_clk;
  wire  readArb_reset;
  wire  readArb_io_in_0_ready;
  wire  readArb_io_in_0_valid;
  wire [3:0] readArb_io_in_0_bits_way_en;
  wire [11:0] readArb_io_in_0_bits_addr;
  wire  readArb_io_in_1_ready;
  wire  readArb_io_in_1_valid;
  wire [3:0] readArb_io_in_1_bits_way_en;
  wire [11:0] readArb_io_in_1_bits_addr;
  wire  readArb_io_in_2_ready;
  wire  readArb_io_in_2_valid;
  wire [3:0] readArb_io_in_2_bits_way_en;
  wire [11:0] readArb_io_in_2_bits_addr;
  wire  readArb_io_in_3_ready;
  wire  readArb_io_in_3_valid;
  wire [3:0] readArb_io_in_3_bits_way_en;
  wire [11:0] readArb_io_in_3_bits_addr;
  wire  readArb_io_out_ready;
  wire  readArb_io_out_valid;
  wire [3:0] readArb_io_out_bits_way_en;
  wire [11:0] readArb_io_out_bits_addr;
  wire [1:0] readArb_io_chosen;
  wire  writeArb_clk;
  wire  writeArb_reset;
  wire  writeArb_io_in_0_ready;
  wire  writeArb_io_in_0_valid;
  wire [3:0] writeArb_io_in_0_bits_way_en;
  wire [11:0] writeArb_io_in_0_bits_addr;
  wire  writeArb_io_in_0_bits_wmask;
  wire [63:0] writeArb_io_in_0_bits_data;
  wire  writeArb_io_in_1_ready;
  wire  writeArb_io_in_1_valid;
  wire [3:0] writeArb_io_in_1_bits_way_en;
  wire [11:0] writeArb_io_in_1_bits_addr;
  wire  writeArb_io_in_1_bits_wmask;
  wire [63:0] writeArb_io_in_1_bits_data;
  wire  writeArb_io_out_ready;
  wire  writeArb_io_out_valid;
  wire [3:0] writeArb_io_out_bits_way_en;
  wire [11:0] writeArb_io_out_bits_addr;
  wire  writeArb_io_out_bits_wmask;
  wire [63:0] writeArb_io_out_bits_data;
  wire  writeArb_io_chosen;
  wire [63:0] T_2770;
  wire [33:0] T_2771;
  wire  T_2773;
  wire  GEN_32;
  wire  T_2778;
  wire  GEN_33;
  wire [33:0] T_2780;
  wire [19:0] T_2783;
  wire  T_2784;
  wire  T_2786;
  wire  T_2788;
  wire  T_2790;
  wire  T_2796_0;
  wire  T_2796_1;
  wire  T_2796_2;
  wire  T_2796_3;
  wire [1:0] T_2798;
  wire [1:0] T_2799;
  wire [3:0] s1_tag_eq_way;
  wire  T_2800;
  wire  T_2801;
  wire  T_2802;
  wire  T_2803;
  wire  T_2804;
  wire  T_2805;
  wire  T_2806;
  wire  T_2807;
  wire  T_2808;
  wire  T_2809;
  wire  T_2810;
  wire  T_2811;
  wire  T_2817_0;
  wire  T_2817_1;
  wire  T_2817_2;
  wire  T_2817_3;
  wire [1:0] T_2819;
  wire [1:0] T_2820;
  wire [3:0] s1_tag_match_way;
  wire  T_2822;
  reg [3:0] s2_tag_match_way;
  reg [31:0] GEN_137;
  wire [3:0] GEN_34;
  wire [3:0] GEN_89;
  wire  s2_tag_match;
  reg [1:0] T_2827_state;
  reg [31:0] GEN_138;
  wire [1:0] GEN_35;
  reg [1:0] T_2852_state;
  reg [31:0] GEN_139;
  wire [1:0] GEN_36;
  reg [1:0] T_2877_state;
  reg [31:0] GEN_140;
  wire [1:0] GEN_37;
  reg [1:0] T_2902_state;
  reg [31:0] GEN_141;
  wire [1:0] GEN_38;
  wire [1:0] T_3124_0_state;
  wire [1:0] T_3124_1_state;
  wire [1:0] T_3124_2_state;
  wire [1:0] T_3124_3_state;
  wire  T_3246;
  wire  T_3247;
  wire  T_3248;
  wire  T_3249;
  wire [1:0] T_3251;
  wire [1:0] T_3253;
  wire [1:0] T_3255;
  wire [1:0] T_3257;
  wire [1:0] T_3283;
  wire [1:0] T_3284;
  wire [1:0] T_3285;
  wire [1:0] s2_hit_state_state;
  wire  T_3336;
  wire  T_3337;
  wire  T_3338;
  wire  T_3339;
  wire  T_3340;
  wire  T_3341;
  wire  T_3342;
  wire  T_3343;
  wire  T_3344;
  wire  T_3345;
  wire  T_3346;
  wire [1:0] T_3352_0;
  wire [1:0] T_3352_1;
  wire  T_3354;
  wire  T_3355;
  wire  T_3358;
  wire [1:0] T_3364_0;
  wire [1:0] T_3364_1;
  wire [1:0] T_3364_2;
  wire  T_3366;
  wire  T_3367;
  wire  T_3368;
  wire  T_3371;
  wire  T_3372;
  wire  T_3373;
  wire  T_3374;
  wire [1:0] T_3382;
  wire [1:0] T_3408_state;
  wire  T_3433;
  wire  s2_hit;
  reg [4:0] lrsc_count;
  reg [31:0] GEN_142;
  wire [4:0] GEN_90;
  wire  lrsc_valid;
  reg [33:0] lrsc_addr;
  reg [63:0] GEN_143;
  wire  T_3438;
  wire  s2_lrsc_addr_match;
  wire  T_3440;
  wire  s2_sc_fail;
  wire [4:0] GEN_91;
  wire [5:0] T_3442;
  wire [4:0] T_3443;
  wire [4:0] GEN_39;
  wire  T_3444;
  wire  T_3445;
  wire  T_3447;
  wire [4:0] GEN_40;
  wire [4:0] GEN_41;
  wire [33:0] GEN_42;
  wire [4:0] GEN_43;
  wire [4:0] GEN_44;
  wire [33:0] GEN_45;
  wire [4:0] GEN_46;
  wire [63:0] s2_data_0;
  wire [63:0] s2_data_1;
  wire [63:0] s2_data_2;
  wire [63:0] s2_data_3;
  reg [63:0] T_3465_0;
  reg [63:0] GEN_144;
  wire  T_3468;
  wire [63:0] T_3476;
  wire [63:0] GEN_47;
  reg [63:0] T_3483_0;
  reg [63:0] GEN_145;
  wire  T_3486;
  wire [63:0] T_3494;
  wire [63:0] GEN_48;
  reg [63:0] T_3501_0;
  reg [63:0] GEN_146;
  wire  T_3504;
  wire [63:0] T_3512;
  wire [63:0] GEN_49;
  reg [63:0] T_3519_0;
  reg [63:0] GEN_147;
  wire  T_3522;
  wire [63:0] T_3530;
  wire [63:0] GEN_50;
  wire [63:0] T_3536;
  wire [63:0] T_3538;
  wire [63:0] T_3540;
  wire [63:0] T_3542;
  wire [63:0] T_3544;
  wire [63:0] T_3545;
  wire [63:0] T_3546;
  wire [63:0] s2_data_muxed;
  wire [63:0] T_3553_0;
  wire [63:0] T_3560_0;
  wire  T_3568_0;
  wire  T_3570;
  wire  T_3574;
  wire  T_3575;
  wire  T_3583;
  wire  amoalu_clk;
  wire  amoalu_reset;
  wire [5:0] amoalu_io_addr;
  wire [4:0] amoalu_io_cmd;
  wire [2:0] amoalu_io_typ;
  wire [63:0] amoalu_io_lhs;
  wire [63:0] amoalu_io_rhs;
  wire [63:0] amoalu_io_out;
  wire  T_3584;
  wire  T_3592;
  wire  T_3593;
  wire [63:0] T_3594;
  wire [39:0] GEN_51;
  wire [8:0] GEN_52;
  wire [4:0] GEN_53;
  wire [2:0] GEN_54;
  wire  GEN_55;
  wire [63:0] GEN_56;
  wire [3:0] GEN_57;
  wire [1:0] GEN_92;
  wire [1:0] rowWMask;
  wire  T_3598;
  reg [15:0] T_3601;
  reg [31:0] GEN_148;
  wire  T_3602;
  wire  T_3603;
  wire  T_3604;
  wire  T_3605;
  wire  T_3606;
  wire  T_3607;
  wire  T_3608;
  wire [14:0] T_3609;
  wire [15:0] T_3610;
  wire [15:0] GEN_58;
  wire [1:0] T_3611;
  wire [3:0] s1_replaced_way_en;
  reg [1:0] T_3614;
  reg [31:0] GEN_149;
  wire [1:0] GEN_59;
  wire [3:0] s2_replaced_way_en;
  wire  T_3616;
  wire  T_3617;
  reg [19:0] T_3618_tag;
  reg [31:0] GEN_150;
  reg [1:0] T_3618_coh_state;
  reg [31:0] GEN_151;
  wire [19:0] GEN_60;
  wire [1:0] GEN_61;
  wire  T_3714;
  wire  T_3715;
  reg [19:0] T_3716_tag;
  reg [31:0] GEN_152;
  reg [1:0] T_3716_coh_state;
  reg [31:0] GEN_153;
  wire [19:0] GEN_62;
  wire [1:0] GEN_63;
  wire  T_3812;
  wire  T_3813;
  reg [19:0] T_3814_tag;
  reg [31:0] GEN_154;
  reg [1:0] T_3814_coh_state;
  reg [31:0] GEN_155;
  wire [19:0] GEN_64;
  wire [1:0] GEN_65;
  wire  T_3910;
  wire  T_3911;
  reg [19:0] T_3912_tag;
  reg [31:0] GEN_156;
  reg [1:0] T_3912_coh_state;
  reg [31:0] GEN_157;
  wire [19:0] GEN_66;
  wire [1:0] GEN_67;
  wire [19:0] T_4773_0_tag;
  wire [1:0] T_4773_0_coh_state;
  wire [19:0] T_4773_1_tag;
  wire [1:0] T_4773_1_coh_state;
  wire [19:0] T_4773_2_tag;
  wire [1:0] T_4773_2_coh_state;
  wire [19:0] T_4773_3_tag;
  wire [1:0] T_4773_3_coh_state;
  wire  T_5250;
  wire  T_5251;
  wire  T_5252;
  wire  T_5253;
  wire [21:0] T_5254;
  wire [21:0] T_5256;
  wire [21:0] T_5257;
  wire [21:0] T_5259;
  wire [21:0] T_5260;
  wire [21:0] T_5262;
  wire [21:0] T_5263;
  wire [21:0] T_5265;
  wire [21:0] T_5362;
  wire [21:0] T_5363;
  wire [21:0] T_5364;
  wire [19:0] s2_repl_meta_tag;
  wire [1:0] s2_repl_meta_coh_state;
  wire [1:0] T_5556;
  wire [19:0] T_5557;
  wire  T_5559;
  wire  T_5560;
  wire  T_5561;
  wire  T_5563;
  wire  T_5564;
  wire  T_5566;
  wire  T_5568;
  wire  T_5572;
  wire  T_5573;
  wire  T_5581;
  wire  T_5582;
  wire [19:0] T_5679_tag;
  wire [1:0] T_5679_coh_state;
  wire [19:0] T_5775_tag;
  wire [1:0] T_5775_coh_state;
  wire [3:0] T_5871;
  wire  T_5872;
  wire  T_5876;
  wire  releaseArb_clk;
  wire  releaseArb_reset;
  wire  releaseArb_io_in_0_ready;
  wire  releaseArb_io_in_0_valid;
  wire [2:0] releaseArb_io_in_0_bits_addr_beat;
  wire [25:0] releaseArb_io_in_0_bits_addr_block;
  wire [1:0] releaseArb_io_in_0_bits_client_xact_id;
  wire  releaseArb_io_in_0_bits_voluntary;
  wire [2:0] releaseArb_io_in_0_bits_r_type;
  wire [63:0] releaseArb_io_in_0_bits_data;
  wire  releaseArb_io_in_1_ready;
  wire  releaseArb_io_in_1_valid;
  wire [2:0] releaseArb_io_in_1_bits_addr_beat;
  wire [25:0] releaseArb_io_in_1_bits_addr_block;
  wire [1:0] releaseArb_io_in_1_bits_client_xact_id;
  wire  releaseArb_io_in_1_bits_voluntary;
  wire [2:0] releaseArb_io_in_1_bits_r_type;
  wire [63:0] releaseArb_io_in_1_bits_data;
  wire  releaseArb_io_out_ready;
  wire  releaseArb_io_out_valid;
  wire [2:0] releaseArb_io_out_bits_addr_beat;
  wire [25:0] releaseArb_io_out_bits_addr_block;
  wire [1:0] releaseArb_io_out_bits_client_xact_id;
  wire  releaseArb_io_out_bits_voluntary;
  wire [2:0] releaseArb_io_out_bits_r_type;
  wire [63:0] releaseArb_io_out_bits_data;
  wire  releaseArb_io_chosen;
  wire  T_5909;
  wire  T_5912;
  wire  FlowThroughSerializer_1_1_clk;
  wire  FlowThroughSerializer_1_1_reset;
  wire  FlowThroughSerializer_1_1_io_in_ready;
  wire  FlowThroughSerializer_1_1_io_in_valid;
  wire [2:0] FlowThroughSerializer_1_1_io_in_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_1_1_io_in_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_1_1_io_in_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_1_io_in_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_1_io_in_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_1_io_in_bits_data;
  wire  FlowThroughSerializer_1_1_io_in_bits_manager_id;
  wire  FlowThroughSerializer_1_1_io_out_ready;
  wire  FlowThroughSerializer_1_1_io_out_valid;
  wire [2:0] FlowThroughSerializer_1_1_io_out_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_1_1_io_out_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_1_1_io_out_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_1_io_out_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_1_io_out_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_1_io_out_bits_data;
  wire  FlowThroughSerializer_1_1_io_out_bits_manager_id;
  wire  FlowThroughSerializer_1_1_io_cnt;
  wire  FlowThroughSerializer_1_1_io_done;
  wire  T_5913;
  wire [2:0] T_5921_0;
  wire [2:0] T_5921_1;
  wire [3:0] GEN_95;
  wire  T_5923;
  wire [3:0] GEN_96;
  wire  T_5924;
  wire  T_5927;
  wire [1:0] T_5933_0;
  wire [1:0] T_5933_1;
  wire [3:0] GEN_97;
  wire  T_5935;
  wire [3:0] GEN_98;
  wire  T_5936;
  wire  T_5939;
  wire  T_5940;
  wire  T_5942;
  wire  T_5943;
  wire [2:0] T_5951_0;
  wire [2:0] T_5951_1;
  wire [3:0] GEN_99;
  wire  T_5953;
  wire [3:0] GEN_100;
  wire  T_5954;
  wire  T_5957;
  wire [1:0] T_5963_0;
  wire [1:0] T_5963_1;
  wire [3:0] GEN_101;
  wire  T_5965;
  wire [3:0] GEN_102;
  wire  T_5966;
  wire  T_5969;
  wire  T_5970;
  wire  T_5971;
  wire  T_5973;
  wire  T_5974;
  wire [63:0] T_5977;
  wire  T_5979;
  wire  T_5980;
  wire  wbArb_clk;
  wire  wbArb_reset;
  wire  wbArb_io_in_0_ready;
  wire  wbArb_io_in_0_valid;
  wire [2:0] wbArb_io_in_0_bits_addr_beat;
  wire [25:0] wbArb_io_in_0_bits_addr_block;
  wire [1:0] wbArb_io_in_0_bits_client_xact_id;
  wire  wbArb_io_in_0_bits_voluntary;
  wire [2:0] wbArb_io_in_0_bits_r_type;
  wire [63:0] wbArb_io_in_0_bits_data;
  wire [3:0] wbArb_io_in_0_bits_way_en;
  wire  wbArb_io_in_1_ready;
  wire  wbArb_io_in_1_valid;
  wire [2:0] wbArb_io_in_1_bits_addr_beat;
  wire [25:0] wbArb_io_in_1_bits_addr_block;
  wire [1:0] wbArb_io_in_1_bits_client_xact_id;
  wire  wbArb_io_in_1_bits_voluntary;
  wire [2:0] wbArb_io_in_1_bits_r_type;
  wire [63:0] wbArb_io_in_1_bits_data;
  wire [3:0] wbArb_io_in_1_bits_way_en;
  wire  wbArb_io_out_ready;
  wire  wbArb_io_out_valid;
  wire [2:0] wbArb_io_out_bits_addr_beat;
  wire [25:0] wbArb_io_out_bits_addr_block;
  wire [1:0] wbArb_io_out_bits_client_xact_id;
  wire  wbArb_io_out_bits_voluntary;
  wire [2:0] wbArb_io_out_bits_r_type;
  wire [63:0] wbArb_io_out_bits_data;
  wire [3:0] wbArb_io_out_bits_way_en;
  wire  wbArb_io_chosen;
  reg  s4_valid;
  reg [31:0] GEN_158;
  wire  T_6036;
  reg [39:0] s4_req_addr;
  reg [63:0] GEN_159;
  reg [8:0] s4_req_tag;
  reg [31:0] GEN_160;
  reg [4:0] s4_req_cmd;
  reg [31:0] GEN_161;
  reg [2:0] s4_req_typ;
  reg [31:0] GEN_162;
  reg  s4_req_phys;
  reg [31:0] GEN_163;
  reg [63:0] s4_req_data;
  reg [63:0] GEN_164;
  wire [39:0] GEN_69;
  wire [8:0] GEN_70;
  wire [4:0] GEN_71;
  wire [2:0] GEN_72;
  wire  GEN_73;
  wire [63:0] GEN_74;
  wire  T_6112;
  wire  T_6115;
  wire [28:0] T_6116;
  wire [36:0] T_6117;
  wire [36:0] GEN_103;
  wire  T_6118;
  wire  T_6119;
  wire  T_6127;
  wire [36:0] T_6129;
  wire  T_6130;
  wire  T_6131;
  wire  T_6132;
  wire  T_6133;
  wire  T_6134;
  wire  T_6135;
  wire  T_6136;
  wire  T_6137;
  wire  T_6138;
  wire  T_6139;
  wire [36:0] T_6141;
  wire  T_6142;
  wire  T_6143;
  wire  T_6144;
  wire  T_6145;
  wire  T_6146;
  wire  T_6147;
  wire  T_6148;
  wire  T_6149;
  wire  T_6150;
  wire  T_6151;
  reg [63:0] s2_store_bypass_data;
  reg [63:0] GEN_165;
  reg  s2_store_bypass;
  reg [31:0] GEN_166;
  wire  T_6155;
  wire  T_6156;
  wire [63:0] T_6157;
  wire [63:0] T_6158;
  wire [63:0] GEN_75;
  wire  GEN_77;
  wire [63:0] GEN_78;
  wire [63:0] s2_data_word_prebypass;
  wire [63:0] s2_data_word;
  wire [1:0] T_6162;
  wire [2:0] T_6163;
  wire  GEN_106;
  wire [2:0] GEN_107;
  wire  T_6165;
  wire  T_6166;
  wire [5:0] T_6167;
  wire  T_6168;
  wire  T_6170;
  wire  T_6171;
  wire  s1_nack;
  wire  T_6172;
  reg  s2_nack_hit;
  reg [31:0] GEN_167;
  wire  GEN_79;
  wire  GEN_80;
  wire  s2_nack_victim;
  wire  T_6177;
  wire  s2_nack_miss;
  wire  T_6178;
  wire  s2_nack;
  wire  T_6180;
  wire  T_6181;
  wire  T_6183;
  wire  s2_recycle_ecc;
  reg  s2_recycle_next;
  reg [31:0] GEN_168;
  wire  GEN_81;
  wire  T_6186;
  reg  block_miss;
  reg [31:0] GEN_169;
  wire  T_6188;
  wire  T_6189;
  wire  GEN_82;
  wire  cache_resp_valid;
  wire [39:0] cache_resp_bits_addr;
  wire [8:0] cache_resp_bits_tag;
  wire [4:0] cache_resp_bits_cmd;
  wire [2:0] cache_resp_bits_typ;
  wire [63:0] cache_resp_bits_data;
  wire  cache_resp_bits_replay;
  wire  cache_resp_bits_has_data;
  wire [63:0] cache_resp_bits_data_word_bypass;
  wire [63:0] cache_resp_bits_store_data;
  wire  T_6590;
  wire  T_6592;
  wire  T_6593;
  wire  T_6603;
  wire [31:0] T_6604;
  wire [31:0] T_6605;
  wire [31:0] T_6606;
  wire  T_6612;
  wire  T_6614;
  wire  T_6615;
  wire [31:0] GEN_108;
  wire [32:0] T_6617;
  wire [31:0] T_6618;
  wire [31:0] T_6620;
  wire [63:0] T_6621;
  wire  T_6622;
  wire [15:0] T_6623;
  wire [15:0] T_6624;
  wire [15:0] T_6625;
  wire  T_6631;
  wire  T_6633;
  wire  T_6634;
  wire [47:0] GEN_110;
  wire [48:0] T_6636;
  wire [47:0] T_6637;
  wire [47:0] T_6638;
  wire [47:0] T_6639;
  wire [63:0] T_6640;
  wire  T_6641;
  wire [7:0] T_6642;
  wire [7:0] T_6643;
  wire [7:0] T_6644;
  wire [7:0] T_6648;
  wire [1:0] GEN_111;
  wire  T_6650;
  wire  T_6651;
  wire  T_6652;
  wire  T_6653;
  wire [55:0] GEN_112;
  wire [56:0] T_6655;
  wire [55:0] T_6656;
  wire [55:0] T_6657;
  wire [55:0] T_6658;
  wire [63:0] T_6659;
  wire [63:0] GEN_113;
  wire [63:0] T_6660;
  wire  uncache_resp_valid;
  wire [39:0] uncache_resp_bits_addr;
  wire [8:0] uncache_resp_bits_tag;
  wire [4:0] uncache_resp_bits_cmd;
  wire [2:0] uncache_resp_bits_typ;
  wire [63:0] uncache_resp_bits_data;
  wire  uncache_resp_bits_replay;
  wire  uncache_resp_bits_has_data;
  wire [63:0] uncache_resp_bits_data_word_bypass;
  wire [63:0] uncache_resp_bits_store_data;
  wire  T_7061;
  reg  T_7062;
  reg [31:0] GEN_170;
  wire  T_7063;
  wire  T_7064_valid;
  wire [39:0] T_7064_bits_addr;
  wire [8:0] T_7064_bits_tag;
  wire [4:0] T_7064_bits_cmd;
  wire [2:0] T_7064_bits_typ;
  wire [63:0] T_7064_bits_data;
  wire  T_7064_bits_replay;
  wire  T_7064_bits_has_data;
  wire [63:0] T_7064_bits_store_data;
  wire  T_7245;
  wire  T_7247;
  wire  T_7248;
  wire  T_7249;
  wire  T_7250;
  reg [1:0] GEN_68;
  reg [31:0] GEN_171;
  reg [3:0] GEN_76;
  reg [31:0] GEN_172;
  reg [3:0] GEN_86;
  reg [31:0] GEN_173;
  reg [63:0] GEN_93;
  reg [63:0] GEN_174;
  WritebackUnit wb (
    .clk(wb_clk),
    .reset(wb_reset),
    .io_req_ready(wb_io_req_ready),
    .io_req_valid(wb_io_req_valid),
    .io_req_bits_addr_beat(wb_io_req_bits_addr_beat),
    .io_req_bits_addr_block(wb_io_req_bits_addr_block),
    .io_req_bits_client_xact_id(wb_io_req_bits_client_xact_id),
    .io_req_bits_voluntary(wb_io_req_bits_voluntary),
    .io_req_bits_r_type(wb_io_req_bits_r_type),
    .io_req_bits_data(wb_io_req_bits_data),
    .io_req_bits_way_en(wb_io_req_bits_way_en),
    .io_meta_read_ready(wb_io_meta_read_ready),
    .io_meta_read_valid(wb_io_meta_read_valid),
    .io_meta_read_bits_idx(wb_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(wb_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(wb_io_meta_read_bits_tag),
    .io_data_req_ready(wb_io_data_req_ready),
    .io_data_req_valid(wb_io_data_req_valid),
    .io_data_req_bits_way_en(wb_io_data_req_bits_way_en),
    .io_data_req_bits_addr(wb_io_data_req_bits_addr),
    .io_data_resp(wb_io_data_resp),
    .io_release_ready(wb_io_release_ready),
    .io_release_valid(wb_io_release_valid),
    .io_release_bits_addr_beat(wb_io_release_bits_addr_beat),
    .io_release_bits_addr_block(wb_io_release_bits_addr_block),
    .io_release_bits_client_xact_id(wb_io_release_bits_client_xact_id),
    .io_release_bits_voluntary(wb_io_release_bits_voluntary),
    .io_release_bits_r_type(wb_io_release_bits_r_type),
    .io_release_bits_data(wb_io_release_bits_data)
  );
  ProbeUnit prober (
    .clk(prober_clk),
    .reset(prober_reset),
    .io_req_ready(prober_io_req_ready),
    .io_req_valid(prober_io_req_valid),
    .io_req_bits_addr_block(prober_io_req_bits_addr_block),
    .io_req_bits_p_type(prober_io_req_bits_p_type),
    .io_req_bits_client_xact_id(prober_io_req_bits_client_xact_id),
    .io_rep_ready(prober_io_rep_ready),
    .io_rep_valid(prober_io_rep_valid),
    .io_rep_bits_addr_beat(prober_io_rep_bits_addr_beat),
    .io_rep_bits_addr_block(prober_io_rep_bits_addr_block),
    .io_rep_bits_client_xact_id(prober_io_rep_bits_client_xact_id),
    .io_rep_bits_voluntary(prober_io_rep_bits_voluntary),
    .io_rep_bits_r_type(prober_io_rep_bits_r_type),
    .io_rep_bits_data(prober_io_rep_bits_data),
    .io_meta_read_ready(prober_io_meta_read_ready),
    .io_meta_read_valid(prober_io_meta_read_valid),
    .io_meta_read_bits_idx(prober_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(prober_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(prober_io_meta_read_bits_tag),
    .io_meta_write_ready(prober_io_meta_write_ready),
    .io_meta_write_valid(prober_io_meta_write_valid),
    .io_meta_write_bits_idx(prober_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(prober_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(prober_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(prober_io_meta_write_bits_data_coh_state),
    .io_wb_req_ready(prober_io_wb_req_ready),
    .io_wb_req_valid(prober_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(prober_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(prober_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(prober_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(prober_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(prober_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(prober_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(prober_io_wb_req_bits_way_en),
    .io_way_en(prober_io_way_en),
    .io_mshr_rdy(prober_io_mshr_rdy),
    .io_block_state_state(prober_io_block_state_state)
  );
  MSHRFile mshrs (
    .clk(mshrs_clk),
    .reset(mshrs_reset),
    .io_req_ready(mshrs_io_req_ready),
    .io_req_valid(mshrs_io_req_valid),
    .io_req_bits_addr(mshrs_io_req_bits_addr),
    .io_req_bits_tag(mshrs_io_req_bits_tag),
    .io_req_bits_cmd(mshrs_io_req_bits_cmd),
    .io_req_bits_typ(mshrs_io_req_bits_typ),
    .io_req_bits_phys(mshrs_io_req_bits_phys),
    .io_req_bits_data(mshrs_io_req_bits_data),
    .io_req_bits_tag_match(mshrs_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(mshrs_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(mshrs_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(mshrs_io_req_bits_way_en),
    .io_resp_ready(mshrs_io_resp_ready),
    .io_resp_valid(mshrs_io_resp_valid),
    .io_resp_bits_addr(mshrs_io_resp_bits_addr),
    .io_resp_bits_tag(mshrs_io_resp_bits_tag),
    .io_resp_bits_cmd(mshrs_io_resp_bits_cmd),
    .io_resp_bits_typ(mshrs_io_resp_bits_typ),
    .io_resp_bits_data(mshrs_io_resp_bits_data),
    .io_resp_bits_replay(mshrs_io_resp_bits_replay),
    .io_resp_bits_has_data(mshrs_io_resp_bits_has_data),
    .io_resp_bits_data_word_bypass(mshrs_io_resp_bits_data_word_bypass),
    .io_resp_bits_store_data(mshrs_io_resp_bits_store_data),
    .io_secondary_miss(mshrs_io_secondary_miss),
    .io_mem_req_ready(mshrs_io_mem_req_ready),
    .io_mem_req_valid(mshrs_io_mem_req_valid),
    .io_mem_req_bits_addr_block(mshrs_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(mshrs_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(mshrs_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(mshrs_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(mshrs_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(mshrs_io_mem_req_bits_union),
    .io_mem_req_bits_data(mshrs_io_mem_req_bits_data),
    .io_refill_way_en(mshrs_io_refill_way_en),
    .io_refill_addr(mshrs_io_refill_addr),
    .io_meta_read_ready(mshrs_io_meta_read_ready),
    .io_meta_read_valid(mshrs_io_meta_read_valid),
    .io_meta_read_bits_idx(mshrs_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(mshrs_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(mshrs_io_meta_read_bits_tag),
    .io_meta_write_ready(mshrs_io_meta_write_ready),
    .io_meta_write_valid(mshrs_io_meta_write_valid),
    .io_meta_write_bits_idx(mshrs_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(mshrs_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(mshrs_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(mshrs_io_meta_write_bits_data_coh_state),
    .io_replay_ready(mshrs_io_replay_ready),
    .io_replay_valid(mshrs_io_replay_valid),
    .io_replay_bits_addr(mshrs_io_replay_bits_addr),
    .io_replay_bits_tag(mshrs_io_replay_bits_tag),
    .io_replay_bits_cmd(mshrs_io_replay_bits_cmd),
    .io_replay_bits_typ(mshrs_io_replay_bits_typ),
    .io_replay_bits_phys(mshrs_io_replay_bits_phys),
    .io_replay_bits_data(mshrs_io_replay_bits_data),
    .io_mem_grant_valid(mshrs_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(mshrs_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(mshrs_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(mshrs_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(mshrs_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(mshrs_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(mshrs_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(mshrs_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(mshrs_io_mem_finish_ready),
    .io_mem_finish_valid(mshrs_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(mshrs_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(mshrs_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(mshrs_io_wb_req_ready),
    .io_wb_req_valid(mshrs_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(mshrs_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(mshrs_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(mshrs_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(mshrs_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(mshrs_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(mshrs_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(mshrs_io_wb_req_bits_way_en),
    .io_probe_rdy(mshrs_io_probe_rdy),
    .io_fence_rdy(mshrs_io_fence_rdy),
    .io_replay_next(mshrs_io_replay_next)
  );
  TLB dtlb (
    .clk(dtlb_clk),
    .reset(dtlb_reset),
    .io_req_ready(dtlb_io_req_ready),
    .io_req_valid(dtlb_io_req_valid),
    .io_req_bits_vpn(dtlb_io_req_bits_vpn),
    .io_req_bits_passthrough(dtlb_io_req_bits_passthrough),
    .io_req_bits_instruction(dtlb_io_req_bits_instruction),
    .io_req_bits_store(dtlb_io_req_bits_store),
    .io_resp_miss(dtlb_io_resp_miss),
    .io_resp_ppn(dtlb_io_resp_ppn),
    .io_resp_xcpt_ld(dtlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(dtlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(dtlb_io_resp_xcpt_if),
    .io_resp_hit_idx(dtlb_io_resp_hit_idx),
    .io_ptw_req_ready(dtlb_io_ptw_req_ready),
    .io_ptw_req_valid(dtlb_io_ptw_req_valid),
    .io_ptw_req_bits_addr(dtlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_prv(dtlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_store(dtlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(dtlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(dtlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_ppn(dtlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(dtlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(dtlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_r(dtlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_typ(dtlb_io_ptw_resp_bits_pte_typ),
    .io_ptw_resp_bits_pte_v(dtlb_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(dtlb_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(dtlb_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(dtlb_io_ptw_invalidate),
    .io_ptw_status_debug(dtlb_io_ptw_status_debug),
    .io_ptw_status_prv(dtlb_io_ptw_status_prv),
    .io_ptw_status_sd(dtlb_io_ptw_status_sd),
    .io_ptw_status_zero3(dtlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(dtlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(dtlb_io_ptw_status_zero2),
    .io_ptw_status_vm(dtlb_io_ptw_status_vm),
    .io_ptw_status_zero1(dtlb_io_ptw_status_zero1),
    .io_ptw_status_pum(dtlb_io_ptw_status_pum),
    .io_ptw_status_mprv(dtlb_io_ptw_status_mprv),
    .io_ptw_status_xs(dtlb_io_ptw_status_xs),
    .io_ptw_status_fs(dtlb_io_ptw_status_fs),
    .io_ptw_status_mpp(dtlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(dtlb_io_ptw_status_hpp),
    .io_ptw_status_spp(dtlb_io_ptw_status_spp),
    .io_ptw_status_mpie(dtlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(dtlb_io_ptw_status_hpie),
    .io_ptw_status_spie(dtlb_io_ptw_status_spie),
    .io_ptw_status_upie(dtlb_io_ptw_status_upie),
    .io_ptw_status_mie(dtlb_io_ptw_status_mie),
    .io_ptw_status_hie(dtlb_io_ptw_status_hie),
    .io_ptw_status_sie(dtlb_io_ptw_status_sie),
    .io_ptw_status_uie(dtlb_io_ptw_status_uie)
  );
  MetadataArray meta (
    .clk(meta_clk),
    .reset(meta_reset),
    .io_read_ready(meta_io_read_ready),
    .io_read_valid(meta_io_read_valid),
    .io_read_bits_idx(meta_io_read_bits_idx),
    .io_read_bits_way_en(meta_io_read_bits_way_en),
    .io_write_ready(meta_io_write_ready),
    .io_write_valid(meta_io_write_valid),
    .io_write_bits_idx(meta_io_write_bits_idx),
    .io_write_bits_way_en(meta_io_write_bits_way_en),
    .io_write_bits_data_tag(meta_io_write_bits_data_tag),
    .io_write_bits_data_coh_state(meta_io_write_bits_data_coh_state),
    .io_resp_0_tag(meta_io_resp_0_tag),
    .io_resp_0_coh_state(meta_io_resp_0_coh_state),
    .io_resp_1_tag(meta_io_resp_1_tag),
    .io_resp_1_coh_state(meta_io_resp_1_coh_state),
    .io_resp_2_tag(meta_io_resp_2_tag),
    .io_resp_2_coh_state(meta_io_resp_2_coh_state),
    .io_resp_3_tag(meta_io_resp_3_tag),
    .io_resp_3_coh_state(meta_io_resp_3_coh_state)
  );
  Arbiter_8 metaReadArb (
    .clk(metaReadArb_clk),
    .reset(metaReadArb_reset),
    .io_in_0_ready(metaReadArb_io_in_0_ready),
    .io_in_0_valid(metaReadArb_io_in_0_valid),
    .io_in_0_bits_idx(metaReadArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaReadArb_io_in_0_bits_way_en),
    .io_in_1_ready(metaReadArb_io_in_1_ready),
    .io_in_1_valid(metaReadArb_io_in_1_valid),
    .io_in_1_bits_idx(metaReadArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaReadArb_io_in_1_bits_way_en),
    .io_in_2_ready(metaReadArb_io_in_2_ready),
    .io_in_2_valid(metaReadArb_io_in_2_valid),
    .io_in_2_bits_idx(metaReadArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaReadArb_io_in_2_bits_way_en),
    .io_in_3_ready(metaReadArb_io_in_3_ready),
    .io_in_3_valid(metaReadArb_io_in_3_valid),
    .io_in_3_bits_idx(metaReadArb_io_in_3_bits_idx),
    .io_in_3_bits_way_en(metaReadArb_io_in_3_bits_way_en),
    .io_in_4_ready(metaReadArb_io_in_4_ready),
    .io_in_4_valid(metaReadArb_io_in_4_valid),
    .io_in_4_bits_idx(metaReadArb_io_in_4_bits_idx),
    .io_in_4_bits_way_en(metaReadArb_io_in_4_bits_way_en),
    .io_out_ready(metaReadArb_io_out_ready),
    .io_out_valid(metaReadArb_io_out_valid),
    .io_out_bits_idx(metaReadArb_io_out_bits_idx),
    .io_out_bits_way_en(metaReadArb_io_out_bits_way_en),
    .io_chosen(metaReadArb_io_chosen)
  );
  Arbiter_1 metaWriteArb (
    .clk(metaWriteArb_clk),
    .reset(metaWriteArb_reset),
    .io_in_0_ready(metaWriteArb_io_in_0_ready),
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_idx(metaWriteArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaWriteArb_io_in_0_bits_way_en),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_coh_state(metaWriteArb_io_in_0_bits_data_coh_state),
    .io_in_1_ready(metaWriteArb_io_in_1_ready),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_idx(metaWriteArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaWriteArb_io_in_1_bits_way_en),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_coh_state(metaWriteArb_io_in_1_bits_data_coh_state),
    .io_out_ready(metaWriteArb_io_out_ready),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_idx(metaWriteArb_io_out_bits_idx),
    .io_out_bits_way_en(metaWriteArb_io_out_bits_way_en),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_coh_state(metaWriteArb_io_out_bits_data_coh_state),
    .io_chosen(metaWriteArb_io_chosen)
  );
  DataArray data (
    .clk(data_clk),
    .reset(data_reset),
    .io_read_ready(data_io_read_ready),
    .io_read_valid(data_io_read_valid),
    .io_read_bits_way_en(data_io_read_bits_way_en),
    .io_read_bits_addr(data_io_read_bits_addr),
    .io_write_ready(data_io_write_ready),
    .io_write_valid(data_io_write_valid),
    .io_write_bits_way_en(data_io_write_bits_way_en),
    .io_write_bits_addr(data_io_write_bits_addr),
    .io_write_bits_wmask(data_io_write_bits_wmask),
    .io_write_bits_data(data_io_write_bits_data),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3)
  );
  Arbiter_10 readArb (
    .clk(readArb_clk),
    .reset(readArb_reset),
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_way_en(readArb_io_in_0_bits_way_en),
    .io_in_0_bits_addr(readArb_io_in_0_bits_addr),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_way_en(readArb_io_in_1_bits_way_en),
    .io_in_1_bits_addr(readArb_io_in_1_bits_addr),
    .io_in_2_ready(readArb_io_in_2_ready),
    .io_in_2_valid(readArb_io_in_2_valid),
    .io_in_2_bits_way_en(readArb_io_in_2_bits_way_en),
    .io_in_2_bits_addr(readArb_io_in_2_bits_addr),
    .io_in_3_ready(readArb_io_in_3_ready),
    .io_in_3_valid(readArb_io_in_3_valid),
    .io_in_3_bits_way_en(readArb_io_in_3_bits_way_en),
    .io_in_3_bits_addr(readArb_io_in_3_bits_addr),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_way_en(readArb_io_out_bits_way_en),
    .io_out_bits_addr(readArb_io_out_bits_addr),
    .io_chosen(readArb_io_chosen)
  );
  Arbiter_11 writeArb (
    .clk(writeArb_clk),
    .reset(writeArb_reset),
    .io_in_0_ready(writeArb_io_in_0_ready),
    .io_in_0_valid(writeArb_io_in_0_valid),
    .io_in_0_bits_way_en(writeArb_io_in_0_bits_way_en),
    .io_in_0_bits_addr(writeArb_io_in_0_bits_addr),
    .io_in_0_bits_wmask(writeArb_io_in_0_bits_wmask),
    .io_in_0_bits_data(writeArb_io_in_0_bits_data),
    .io_in_1_ready(writeArb_io_in_1_ready),
    .io_in_1_valid(writeArb_io_in_1_valid),
    .io_in_1_bits_way_en(writeArb_io_in_1_bits_way_en),
    .io_in_1_bits_addr(writeArb_io_in_1_bits_addr),
    .io_in_1_bits_wmask(writeArb_io_in_1_bits_wmask),
    .io_in_1_bits_data(writeArb_io_in_1_bits_data),
    .io_out_ready(writeArb_io_out_ready),
    .io_out_valid(writeArb_io_out_valid),
    .io_out_bits_way_en(writeArb_io_out_bits_way_en),
    .io_out_bits_addr(writeArb_io_out_bits_addr),
    .io_out_bits_wmask(writeArb_io_out_bits_wmask),
    .io_out_bits_data(writeArb_io_out_bits_data),
    .io_chosen(writeArb_io_chosen)
  );
  AMOALU amoalu (
    .clk(amoalu_clk),
    .reset(amoalu_reset),
    .io_addr(amoalu_io_addr),
    .io_cmd(amoalu_io_cmd),
    .io_typ(amoalu_io_typ),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out)
  );
  LockingArbiter_1 releaseArb (
    .clk(releaseArb_clk),
    .reset(releaseArb_reset),
    .io_in_0_ready(releaseArb_io_in_0_ready),
    .io_in_0_valid(releaseArb_io_in_0_valid),
    .io_in_0_bits_addr_beat(releaseArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(releaseArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(releaseArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(releaseArb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(releaseArb_io_in_0_bits_r_type),
    .io_in_0_bits_data(releaseArb_io_in_0_bits_data),
    .io_in_1_ready(releaseArb_io_in_1_ready),
    .io_in_1_valid(releaseArb_io_in_1_valid),
    .io_in_1_bits_addr_beat(releaseArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(releaseArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(releaseArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(releaseArb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(releaseArb_io_in_1_bits_r_type),
    .io_in_1_bits_data(releaseArb_io_in_1_bits_data),
    .io_out_ready(releaseArb_io_out_ready),
    .io_out_valid(releaseArb_io_out_valid),
    .io_out_bits_addr_beat(releaseArb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(releaseArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(releaseArb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(releaseArb_io_out_bits_voluntary),
    .io_out_bits_r_type(releaseArb_io_out_bits_r_type),
    .io_out_bits_data(releaseArb_io_out_bits_data),
    .io_chosen(releaseArb_io_chosen)
  );
  FlowThroughSerializer_1 FlowThroughSerializer_1_1 (
    .clk(FlowThroughSerializer_1_1_clk),
    .reset(FlowThroughSerializer_1_1_reset),
    .io_in_ready(FlowThroughSerializer_1_1_io_in_ready),
    .io_in_valid(FlowThroughSerializer_1_1_io_in_valid),
    .io_in_bits_addr_beat(FlowThroughSerializer_1_1_io_in_bits_addr_beat),
    .io_in_bits_client_xact_id(FlowThroughSerializer_1_1_io_in_bits_client_xact_id),
    .io_in_bits_manager_xact_id(FlowThroughSerializer_1_1_io_in_bits_manager_xact_id),
    .io_in_bits_is_builtin_type(FlowThroughSerializer_1_1_io_in_bits_is_builtin_type),
    .io_in_bits_g_type(FlowThroughSerializer_1_1_io_in_bits_g_type),
    .io_in_bits_data(FlowThroughSerializer_1_1_io_in_bits_data),
    .io_in_bits_manager_id(FlowThroughSerializer_1_1_io_in_bits_manager_id),
    .io_out_ready(FlowThroughSerializer_1_1_io_out_ready),
    .io_out_valid(FlowThroughSerializer_1_1_io_out_valid),
    .io_out_bits_addr_beat(FlowThroughSerializer_1_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(FlowThroughSerializer_1_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(FlowThroughSerializer_1_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(FlowThroughSerializer_1_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(FlowThroughSerializer_1_1_io_out_bits_g_type),
    .io_out_bits_data(FlowThroughSerializer_1_1_io_out_bits_data),
    .io_out_bits_manager_id(FlowThroughSerializer_1_1_io_out_bits_manager_id),
    .io_cnt(FlowThroughSerializer_1_1_io_cnt),
    .io_done(FlowThroughSerializer_1_1_io_done)
  );
  Arbiter_3 wbArb (
    .clk(wbArb_clk),
    .reset(wbArb_reset),
    .io_in_0_ready(wbArb_io_in_0_ready),
    .io_in_0_valid(wbArb_io_in_0_valid),
    .io_in_0_bits_addr_beat(wbArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(wbArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(wbArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(wbArb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(wbArb_io_in_0_bits_r_type),
    .io_in_0_bits_data(wbArb_io_in_0_bits_data),
    .io_in_0_bits_way_en(wbArb_io_in_0_bits_way_en),
    .io_in_1_ready(wbArb_io_in_1_ready),
    .io_in_1_valid(wbArb_io_in_1_valid),
    .io_in_1_bits_addr_beat(wbArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(wbArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(wbArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(wbArb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(wbArb_io_in_1_bits_r_type),
    .io_in_1_bits_data(wbArb_io_in_1_bits_data),
    .io_in_1_bits_way_en(wbArb_io_in_1_bits_way_en),
    .io_out_ready(wbArb_io_out_ready),
    .io_out_valid(wbArb_io_out_valid),
    .io_out_bits_addr_beat(wbArb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(wbArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(wbArb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(wbArb_io_out_bits_voluntary),
    .io_out_bits_r_type(wbArb_io_out_bits_r_type),
    .io_out_bits_data(wbArb_io_out_bits_data),
    .io_out_bits_way_en(wbArb_io_out_bits_way_en),
    .io_chosen(wbArb_io_chosen)
  );
  assign io_cpu_req_ready = GEN_82;
  assign io_cpu_s2_nack = T_7063;
  assign io_cpu_resp_valid = T_7064_valid;
  assign io_cpu_resp_bits_addr = T_7064_bits_addr;
  assign io_cpu_resp_bits_tag = T_7064_bits_tag;
  assign io_cpu_resp_bits_cmd = T_7064_bits_cmd;
  assign io_cpu_resp_bits_typ = T_7064_bits_typ;
  assign io_cpu_resp_bits_data = T_7064_bits_data;
  assign io_cpu_resp_bits_replay = T_7064_bits_replay;
  assign io_cpu_resp_bits_has_data = T_7064_bits_has_data;
  assign io_cpu_resp_bits_data_word_bypass = T_6621;
  assign io_cpu_resp_bits_store_data = T_7064_bits_store_data;
  assign io_cpu_replay_next = T_7250;
  assign io_cpu_xcpt_ma_ld = T_2366;
  assign io_cpu_xcpt_ma_st = T_2367;
  assign io_cpu_xcpt_pf_ld = T_2368;
  assign io_cpu_xcpt_pf_st = T_2369;
  assign io_cpu_ordered = T_7248;
  assign io_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_ptw_req_bits_addr = dtlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_prv = dtlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_store = dtlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = dtlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = mshrs_io_mem_req_valid;
  assign io_mem_acquire_bits_addr_block = mshrs_io_mem_req_bits_addr_block;
  assign io_mem_acquire_bits_client_xact_id = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = mshrs_io_mem_req_bits_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = mshrs_io_mem_req_bits_is_builtin_type;
  assign io_mem_acquire_bits_a_type = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_union = mshrs_io_mem_req_bits_union;
  assign io_mem_acquire_bits_data = mshrs_io_mem_req_bits_data;
  assign io_mem_probe_ready = T_5912;
  assign io_mem_release_valid = releaseArb_io_out_valid;
  assign io_mem_release_bits_addr_beat = releaseArb_io_out_bits_addr_beat;
  assign io_mem_release_bits_addr_block = releaseArb_io_out_bits_addr_block;
  assign io_mem_release_bits_client_xact_id = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_voluntary = releaseArb_io_out_bits_voluntary;
  assign io_mem_release_bits_r_type = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_data = releaseArb_io_out_bits_data;
  assign io_mem_grant_ready = FlowThroughSerializer_1_1_io_in_ready;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_finish_bits_manager_xact_id = mshrs_io_mem_finish_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = mshrs_io_mem_finish_bits_manager_id;
  assign wb_clk = clk;
  assign wb_reset = reset;
  assign wb_io_req_valid = wbArb_io_out_valid;
  assign wb_io_req_bits_addr_beat = wbArb_io_out_bits_addr_beat;
  assign wb_io_req_bits_addr_block = wbArb_io_out_bits_addr_block;
  assign wb_io_req_bits_client_xact_id = wbArb_io_out_bits_client_xact_id;
  assign wb_io_req_bits_voluntary = wbArb_io_out_bits_voluntary;
  assign wb_io_req_bits_r_type = wbArb_io_out_bits_r_type;
  assign wb_io_req_bits_data = wbArb_io_out_bits_data;
  assign wb_io_req_bits_way_en = wbArb_io_out_bits_way_en;
  assign wb_io_meta_read_ready = metaReadArb_io_in_3_ready;
  assign wb_io_data_req_ready = readArb_io_in_2_ready;
  assign wb_io_data_resp = T_3553_0;
  assign wb_io_release_ready = releaseArb_io_in_0_ready;
  assign prober_clk = clk;
  assign prober_reset = reset;
  assign prober_io_req_valid = T_5909;
  assign prober_io_req_bits_addr_block = io_mem_probe_bits_addr_block;
  assign prober_io_req_bits_p_type = io_mem_probe_bits_p_type;
  assign prober_io_req_bits_client_xact_id = GEN_68;
  assign prober_io_rep_ready = releaseArb_io_in_1_ready;
  assign prober_io_meta_read_ready = metaReadArb_io_in_2_ready;
  assign prober_io_meta_write_ready = metaWriteArb_io_in_1_ready;
  assign prober_io_wb_req_ready = wbArb_io_in_0_ready;
  assign prober_io_way_en = s2_tag_match_way;
  assign prober_io_mshr_rdy = mshrs_io_probe_rdy;
  assign prober_io_block_state_state = s2_hit_state_state;
  assign mshrs_clk = clk;
  assign mshrs_reset = reset;
  assign mshrs_io_req_valid = GEN_80;
  assign mshrs_io_req_bits_addr = s2_req_addr;
  assign mshrs_io_req_bits_tag = s2_req_tag;
  assign mshrs_io_req_bits_cmd = s2_req_cmd;
  assign mshrs_io_req_bits_typ = s2_req_typ;
  assign mshrs_io_req_bits_phys = s2_req_phys;
  assign mshrs_io_req_bits_data = s2_req_data;
  assign mshrs_io_req_bits_tag_match = s2_tag_match;
  assign mshrs_io_req_bits_old_meta_tag = T_5775_tag;
  assign mshrs_io_req_bits_old_meta_coh_state = T_5775_coh_state;
  assign mshrs_io_req_bits_way_en = T_5871;
  assign mshrs_io_resp_ready = T_7062;
  assign mshrs_io_mem_req_ready = io_mem_acquire_ready;
  assign mshrs_io_meta_read_ready = metaReadArb_io_in_1_ready;
  assign mshrs_io_meta_write_ready = metaWriteArb_io_in_0_ready;
  assign mshrs_io_replay_ready = readArb_io_in_1_ready;
  assign mshrs_io_mem_grant_valid = T_5913;
  assign mshrs_io_mem_grant_bits_addr_beat = FlowThroughSerializer_1_1_io_out_bits_addr_beat;
  assign mshrs_io_mem_grant_bits_client_xact_id = FlowThroughSerializer_1_1_io_out_bits_client_xact_id;
  assign mshrs_io_mem_grant_bits_manager_xact_id = FlowThroughSerializer_1_1_io_out_bits_manager_xact_id;
  assign mshrs_io_mem_grant_bits_is_builtin_type = FlowThroughSerializer_1_1_io_out_bits_is_builtin_type;
  assign mshrs_io_mem_grant_bits_g_type = FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign mshrs_io_mem_grant_bits_data = FlowThroughSerializer_1_1_io_out_bits_data;
  assign mshrs_io_mem_grant_bits_manager_id = FlowThroughSerializer_1_1_io_out_bits_manager_id;
  assign mshrs_io_mem_finish_ready = io_mem_finish_ready;
  assign mshrs_io_wb_req_ready = wbArb_io_in_1_ready;
  assign T_2081 = io_cpu_req_ready & io_cpu_req_valid;
  assign T_2159 = io_cpu_s1_kill == 1'h0;
  assign s1_valid_masked = s1_valid & T_2159;
  assign T_2240 = s2_req_cmd != 5'h5;
  assign s2_replay = T_2239 & T_2240;
  assign s2_recycle = T_6186;
  assign s2_valid_masked = T_6181;
  assign GEN_0 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T_2321 = s1_req_cmd == 5'h0;
  assign T_2322 = s1_req_cmd == 5'h6;
  assign T_2323 = T_2321 | T_2322;
  assign T_2324 = s1_req_cmd == 5'h7;
  assign T_2325 = T_2323 | T_2324;
  assign T_2326 = s1_req_cmd[3];
  assign T_2327 = s1_req_cmd == 5'h4;
  assign T_2328 = T_2326 | T_2327;
  assign s1_read = T_2325 | T_2328;
  assign T_2329 = s1_req_cmd == 5'h1;
  assign T_2331 = T_2329 | T_2324;
  assign s1_write = T_2331 | T_2328;
  assign T_2335 = s1_read | s1_write;
  assign T_2336 = s1_req_cmd == 5'h2;
  assign T_2337 = s1_req_cmd == 5'h3;
  assign T_2338 = T_2336 | T_2337;
  assign s1_readwrite = T_2335 | T_2338;
  assign dtlb_clk = clk;
  assign dtlb_reset = reset;
  assign dtlb_io_req_valid = T_2339;
  assign dtlb_io_req_bits_vpn = T_2340;
  assign dtlb_io_req_bits_passthrough = s1_req_phys;
  assign dtlb_io_req_bits_instruction = 1'h0;
  assign dtlb_io_req_bits_store = s1_write;
  assign dtlb_io_ptw_req_ready = io_ptw_req_ready;
  assign dtlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign dtlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign dtlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign dtlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign dtlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign dtlb_io_ptw_resp_bits_pte_typ = io_ptw_resp_bits_pte_typ;
  assign dtlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign dtlb_io_ptw_ptbr_asid = io_ptw_ptbr_asid;
  assign dtlb_io_ptw_ptbr_ppn = io_ptw_ptbr_ppn;
  assign dtlb_io_ptw_invalidate = io_ptw_invalidate;
  assign dtlb_io_ptw_status_debug = io_ptw_status_debug;
  assign dtlb_io_ptw_status_prv = io_ptw_status_prv;
  assign dtlb_io_ptw_status_sd = io_ptw_status_sd;
  assign dtlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign dtlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign dtlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign dtlb_io_ptw_status_vm = io_ptw_status_vm;
  assign dtlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign dtlb_io_ptw_status_pum = io_ptw_status_pum;
  assign dtlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign dtlb_io_ptw_status_xs = io_ptw_status_xs;
  assign dtlb_io_ptw_status_fs = io_ptw_status_fs;
  assign dtlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign dtlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign dtlb_io_ptw_status_spp = io_ptw_status_spp;
  assign dtlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign dtlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign dtlb_io_ptw_status_spie = io_ptw_status_spie;
  assign dtlb_io_ptw_status_upie = io_ptw_status_upie;
  assign dtlb_io_ptw_status_mie = io_ptw_status_mie;
  assign dtlb_io_ptw_status_hie = io_ptw_status_hie;
  assign dtlb_io_ptw_status_sie = io_ptw_status_sie;
  assign dtlb_io_ptw_status_uie = io_ptw_status_uie;
  assign T_2339 = s1_valid_masked & s1_readwrite;
  assign T_2340 = s1_req_addr[39:12];
  assign T_2343 = dtlb_io_req_ready == 1'h0;
  assign T_2345 = io_cpu_req_bits_phys == 1'h0;
  assign T_2346 = T_2343 & T_2345;
  assign GEN_1 = T_2346 ? 1'h0 : 1'h1;
  assign GEN_2 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign GEN_3 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign GEN_4 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign GEN_5 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign GEN_6 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign GEN_7 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T_2348 = {wb_io_meta_read_bits_tag,wb_io_meta_read_bits_idx};
  assign GEN_83 = {{6'd0}, T_2348};
  assign T_2349 = GEN_83 << 6;
  assign GEN_8 = wb_io_meta_read_valid ? {{8'd0}, T_2349} : GEN_2;
  assign GEN_9 = wb_io_meta_read_valid ? 1'h1 : GEN_6;
  assign T_2351 = {prober_io_meta_read_bits_tag,prober_io_meta_read_bits_idx};
  assign GEN_84 = {{6'd0}, T_2351};
  assign T_2352 = GEN_84 << 6;
  assign GEN_10 = prober_io_meta_read_valid ? {{8'd0}, T_2352} : GEN_8;
  assign GEN_11 = prober_io_meta_read_valid ? 1'h1 : GEN_9;
  assign GEN_12 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : GEN_10;
  assign GEN_13 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : GEN_3;
  assign GEN_14 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : GEN_4;
  assign GEN_15 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : GEN_5;
  assign GEN_16 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : GEN_11;
  assign GEN_17 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : GEN_7;
  assign GEN_18 = s2_recycle ? s2_req_addr : GEN_12;
  assign GEN_19 = s2_recycle ? s2_req_tag : GEN_13;
  assign GEN_20 = s2_recycle ? s2_req_cmd : GEN_14;
  assign GEN_21 = s2_recycle ? s2_req_typ : GEN_15;
  assign GEN_22 = s2_recycle ? s2_req_phys : GEN_16;
  assign GEN_23 = s2_recycle ? s2_req_data : GEN_17;
  assign T_2354 = s1_req_addr[11:0];
  assign s1_addr = {dtlb_io_resp_ppn,T_2354};
  assign T_2355 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_s1_data;
  assign GEN_24 = s1_write ? T_2355 : s2_req_data;
  assign GEN_25 = s1_recycled ? s1_req_data : GEN_24;
  assign GEN_26 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign GEN_27 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign GEN_28 = s1_clk_en ? {{8'd0}, s1_addr} : s2_req_addr;
  assign GEN_29 = s1_clk_en ? GEN_25 : s2_req_data;
  assign GEN_30 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign GEN_31 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign T_2357 = s1_req_typ[1:0];
  assign GEN_85 = {{3'd0}, 1'h1};
  assign T_2359 = GEN_85 << T_2357;
  assign T_2361 = T_2359 - GEN_85;
  assign T_2362 = T_2361[3:0];
  assign T_2363 = T_2362[2:0];
  assign GEN_87 = {{37'd0}, T_2363};
  assign T_2364 = s1_req_addr & GEN_87;
  assign GEN_88 = {{39'd0}, 1'h0};
  assign misaligned = T_2364 != GEN_88;
  assign T_2366 = s1_read & misaligned;
  assign T_2367 = s1_write & misaligned;
  assign T_2368 = s1_read & dtlb_io_resp_xcpt_ld;
  assign T_2369 = s1_write & dtlb_io_resp_xcpt_st;
  assign T_2370 = io_cpu_xcpt_ma_ld | io_cpu_xcpt_ma_st;
  assign T_2371 = T_2370 | io_cpu_xcpt_pf_ld;
  assign T_2372 = T_2371 | io_cpu_xcpt_pf_st;
  assign T_2374 = T_2373 & s2_valid_masked;
  assign T_2376 = T_2374 == 1'h0;
  assign T_2377 = T_2376 | reset;
  assign T_2379 = T_2377 == 1'h0;
  assign meta_clk = clk;
  assign meta_reset = reset;
  assign meta_io_read_valid = metaReadArb_io_out_valid;
  assign meta_io_read_bits_idx = metaReadArb_io_out_bits_idx;
  assign meta_io_read_bits_way_en = metaReadArb_io_out_bits_way_en;
  assign meta_io_write_valid = metaWriteArb_io_out_valid;
  assign meta_io_write_bits_idx = metaWriteArb_io_out_bits_idx;
  assign meta_io_write_bits_way_en = metaWriteArb_io_out_bits_way_en;
  assign meta_io_write_bits_data_tag = metaWriteArb_io_out_bits_data_tag;
  assign meta_io_write_bits_data_coh_state = metaWriteArb_io_out_bits_data_coh_state;
  assign metaReadArb_clk = clk;
  assign metaReadArb_reset = reset;
  assign metaReadArb_io_in_0_valid = s2_recycle;
  assign metaReadArb_io_in_0_bits_idx = T_2780[5:0];
  assign metaReadArb_io_in_0_bits_way_en = GEN_76;
  assign metaReadArb_io_in_1_valid = mshrs_io_meta_read_valid;
  assign metaReadArb_io_in_1_bits_idx = mshrs_io_meta_read_bits_idx;
  assign metaReadArb_io_in_1_bits_way_en = mshrs_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_2_valid = prober_io_meta_read_valid;
  assign metaReadArb_io_in_2_bits_idx = prober_io_meta_read_bits_idx;
  assign metaReadArb_io_in_2_bits_way_en = prober_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_3_valid = wb_io_meta_read_valid;
  assign metaReadArb_io_in_3_bits_idx = wb_io_meta_read_bits_idx;
  assign metaReadArb_io_in_3_bits_way_en = wb_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_4_valid = io_cpu_req_valid;
  assign metaReadArb_io_in_4_bits_idx = T_2771[5:0];
  assign metaReadArb_io_in_4_bits_way_en = GEN_86;
  assign metaReadArb_io_out_ready = meta_io_read_ready;
  assign metaWriteArb_clk = clk;
  assign metaWriteArb_reset = reset;
  assign metaWriteArb_io_in_0_valid = mshrs_io_meta_write_valid;
  assign metaWriteArb_io_in_0_bits_idx = mshrs_io_meta_write_bits_idx;
  assign metaWriteArb_io_in_0_bits_way_en = mshrs_io_meta_write_bits_way_en;
  assign metaWriteArb_io_in_0_bits_data_tag = mshrs_io_meta_write_bits_data_tag;
  assign metaWriteArb_io_in_0_bits_data_coh_state = mshrs_io_meta_write_bits_data_coh_state;
  assign metaWriteArb_io_in_1_valid = prober_io_meta_write_valid;
  assign metaWriteArb_io_in_1_bits_idx = prober_io_meta_write_bits_idx;
  assign metaWriteArb_io_in_1_bits_way_en = prober_io_meta_write_bits_way_en;
  assign metaWriteArb_io_in_1_bits_data_tag = prober_io_meta_write_bits_data_tag;
  assign metaWriteArb_io_in_1_bits_data_coh_state = prober_io_meta_write_bits_data_coh_state;
  assign metaWriteArb_io_out_ready = meta_io_write_ready;
  assign data_clk = clk;
  assign data_reset = reset;
  assign data_io_read_valid = readArb_io_out_valid;
  assign data_io_read_bits_way_en = readArb_io_out_bits_way_en;
  assign data_io_read_bits_addr = readArb_io_out_bits_addr;
  assign data_io_write_valid = writeArb_io_out_valid;
  assign data_io_write_bits_way_en = writeArb_io_out_bits_way_en;
  assign data_io_write_bits_addr = writeArb_io_out_bits_addr;
  assign data_io_write_bits_wmask = writeArb_io_out_bits_wmask;
  assign data_io_write_bits_data = T_2770;
  assign readArb_clk = clk;
  assign readArb_reset = reset;
  assign readArb_io_in_0_valid = s2_recycle;
  assign readArb_io_in_0_bits_way_en = 4'hf;
  assign readArb_io_in_0_bits_addr = s2_req_addr[11:0];
  assign readArb_io_in_1_valid = mshrs_io_replay_valid;
  assign readArb_io_in_1_bits_way_en = 4'hf;
  assign readArb_io_in_1_bits_addr = mshrs_io_replay_bits_addr[11:0];
  assign readArb_io_in_2_valid = wb_io_data_req_valid;
  assign readArb_io_in_2_bits_way_en = wb_io_data_req_bits_way_en;
  assign readArb_io_in_2_bits_addr = wb_io_data_req_bits_addr;
  assign readArb_io_in_3_valid = io_cpu_req_valid;
  assign readArb_io_in_3_bits_way_en = 4'hf;
  assign readArb_io_in_3_bits_addr = io_cpu_req_bits_addr[11:0];
  assign readArb_io_out_ready = T_5980;
  assign writeArb_clk = clk;
  assign writeArb_reset = reset;
  assign writeArb_io_in_0_valid = s3_valid;
  assign writeArb_io_in_0_bits_way_en = s3_way;
  assign writeArb_io_in_0_bits_addr = s3_req_addr[11:0];
  assign writeArb_io_in_0_bits_wmask = rowWMask[0];
  assign writeArb_io_in_0_bits_data = s3_req_data;
  assign writeArb_io_in_1_valid = T_5974;
  assign writeArb_io_in_1_bits_way_en = mshrs_io_refill_way_en;
  assign writeArb_io_in_1_bits_addr = mshrs_io_refill_addr;
  assign writeArb_io_in_1_bits_wmask = 1'h1;
  assign writeArb_io_in_1_bits_data = T_5977;
  assign writeArb_io_out_ready = data_io_write_ready;
  assign T_2770 = writeArb_io_out_bits_data;
  assign T_2771 = io_cpu_req_bits_addr[39:6];
  assign T_2773 = metaReadArb_io_in_4_ready == 1'h0;
  assign GEN_32 = T_2773 ? 1'h0 : GEN_1;
  assign T_2778 = readArb_io_in_3_ready == 1'h0;
  assign GEN_33 = T_2778 ? 1'h0 : GEN_32;
  assign T_2780 = s2_req_addr[39:6];
  assign T_2783 = s1_addr[31:12];
  assign T_2784 = meta_io_resp_0_tag == T_2783;
  assign T_2786 = meta_io_resp_1_tag == T_2783;
  assign T_2788 = meta_io_resp_2_tag == T_2783;
  assign T_2790 = meta_io_resp_3_tag == T_2783;
  assign T_2796_0 = T_2784;
  assign T_2796_1 = T_2786;
  assign T_2796_2 = T_2788;
  assign T_2796_3 = T_2790;
  assign T_2798 = {T_2796_1,T_2796_0};
  assign T_2799 = {T_2796_3,T_2796_2};
  assign s1_tag_eq_way = {T_2799,T_2798};
  assign T_2800 = s1_tag_eq_way[0];
  assign T_2801 = meta_io_resp_0_coh_state != 2'h0;
  assign T_2802 = T_2800 & T_2801;
  assign T_2803 = s1_tag_eq_way[1];
  assign T_2804 = meta_io_resp_1_coh_state != 2'h0;
  assign T_2805 = T_2803 & T_2804;
  assign T_2806 = s1_tag_eq_way[2];
  assign T_2807 = meta_io_resp_2_coh_state != 2'h0;
  assign T_2808 = T_2806 & T_2807;
  assign T_2809 = s1_tag_eq_way[3];
  assign T_2810 = meta_io_resp_3_coh_state != 2'h0;
  assign T_2811 = T_2809 & T_2810;
  assign T_2817_0 = T_2802;
  assign T_2817_1 = T_2805;
  assign T_2817_2 = T_2808;
  assign T_2817_3 = T_2811;
  assign T_2819 = {T_2817_1,T_2817_0};
  assign T_2820 = {T_2817_3,T_2817_2};
  assign s1_tag_match_way = {T_2820,T_2819};
  assign T_2822 = s1_valid == 1'h0;
  assign GEN_34 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign GEN_89 = {{3'd0}, 1'h0};
  assign s2_tag_match = s2_tag_match_way != GEN_89;
  assign GEN_35 = s1_clk_en ? meta_io_resp_0_coh_state : T_2827_state;
  assign GEN_36 = s1_clk_en ? meta_io_resp_1_coh_state : T_2852_state;
  assign GEN_37 = s1_clk_en ? meta_io_resp_2_coh_state : T_2877_state;
  assign GEN_38 = s1_clk_en ? meta_io_resp_3_coh_state : T_2902_state;
  assign T_3124_0_state = T_2827_state;
  assign T_3124_1_state = T_2852_state;
  assign T_3124_2_state = T_2877_state;
  assign T_3124_3_state = T_2902_state;
  assign T_3246 = s2_tag_match_way[0];
  assign T_3247 = s2_tag_match_way[1];
  assign T_3248 = s2_tag_match_way[2];
  assign T_3249 = s2_tag_match_way[3];
  assign T_3251 = T_3246 ? T_3124_0_state : {{1'd0}, 1'h0};
  assign T_3253 = T_3247 ? T_3124_1_state : {{1'd0}, 1'h0};
  assign T_3255 = T_3248 ? T_3124_2_state : {{1'd0}, 1'h0};
  assign T_3257 = T_3249 ? T_3124_3_state : {{1'd0}, 1'h0};
  assign T_3283 = T_3251 | T_3253;
  assign T_3284 = T_3283 | T_3255;
  assign T_3285 = T_3284 | T_3257;
  assign s2_hit_state_state = T_3285;
  assign T_3336 = s2_req_cmd == 5'h1;
  assign T_3337 = s2_req_cmd == 5'h7;
  assign T_3338 = T_3336 | T_3337;
  assign T_3339 = s2_req_cmd[3];
  assign T_3340 = s2_req_cmd == 5'h4;
  assign T_3341 = T_3339 | T_3340;
  assign T_3342 = T_3338 | T_3341;
  assign T_3343 = s2_req_cmd == 5'h3;
  assign T_3344 = T_3342 | T_3343;
  assign T_3345 = s2_req_cmd == 5'h6;
  assign T_3346 = T_3344 | T_3345;
  assign T_3352_0 = 2'h2;
  assign T_3352_1 = 2'h3;
  assign T_3354 = T_3352_0 == s2_hit_state_state;
  assign T_3355 = T_3352_1 == s2_hit_state_state;
  assign T_3358 = T_3354 | T_3355;
  assign T_3364_0 = 2'h1;
  assign T_3364_1 = 2'h2;
  assign T_3364_2 = 2'h3;
  assign T_3366 = T_3364_0 == s2_hit_state_state;
  assign T_3367 = T_3364_1 == s2_hit_state_state;
  assign T_3368 = T_3364_2 == s2_hit_state_state;
  assign T_3371 = T_3366 | T_3367;
  assign T_3372 = T_3371 | T_3368;
  assign T_3373 = T_3346 ? T_3358 : T_3372;
  assign T_3374 = s2_tag_match & T_3373;
  assign T_3382 = T_3342 ? 2'h3 : s2_hit_state_state;
  assign T_3408_state = T_3382;
  assign T_3433 = s2_hit_state_state == T_3408_state;
  assign s2_hit = T_3374 & T_3433;
  assign GEN_90 = {{4'd0}, 1'h0};
  assign lrsc_valid = lrsc_count != GEN_90;
  assign T_3438 = lrsc_addr == T_2780;
  assign s2_lrsc_addr_match = lrsc_valid & T_3438;
  assign T_3440 = s2_lrsc_addr_match == 1'h0;
  assign s2_sc_fail = T_3337 & T_3440;
  assign GEN_91 = {{4'd0}, 1'h1};
  assign T_3442 = lrsc_count - GEN_91;
  assign T_3443 = T_3442[4:0];
  assign GEN_39 = lrsc_valid ? T_3443 : lrsc_count;
  assign T_3444 = s2_valid_masked & s2_hit;
  assign T_3445 = T_3444 | s2_replay;
  assign T_3447 = lrsc_valid == 1'h0;
  assign GEN_40 = T_3447 ? 5'h1f : GEN_39;
  assign GEN_41 = T_3345 ? GEN_40 : GEN_39;
  assign GEN_42 = T_3345 ? T_2780 : lrsc_addr;
  assign GEN_43 = T_3337 ? {{4'd0}, 1'h0} : GEN_41;
  assign GEN_44 = T_3445 ? GEN_43 : GEN_39;
  assign GEN_45 = T_3445 ? GEN_42 : lrsc_addr;
  assign GEN_46 = io_cpu_invalidate_lr ? {{4'd0}, 1'h0} : GEN_44;
  assign s2_data_0 = T_3465_0;
  assign s2_data_1 = T_3483_0;
  assign s2_data_2 = T_3501_0;
  assign s2_data_3 = T_3519_0;
  assign T_3468 = s1_clk_en & T_2800;
  assign T_3476 = data_io_resp_0;
  assign GEN_47 = T_3468 ? T_3476 : T_3465_0;
  assign T_3486 = s1_clk_en & T_2803;
  assign T_3494 = data_io_resp_1;
  assign GEN_48 = T_3486 ? T_3494 : T_3483_0;
  assign T_3504 = s1_clk_en & T_2806;
  assign T_3512 = data_io_resp_2;
  assign GEN_49 = T_3504 ? T_3512 : T_3501_0;
  assign T_3522 = s1_clk_en & T_2809;
  assign T_3530 = data_io_resp_3;
  assign GEN_50 = T_3522 ? T_3530 : T_3519_0;
  assign T_3536 = T_3246 ? s2_data_0 : {{63'd0}, 1'h0};
  assign T_3538 = T_3247 ? s2_data_1 : {{63'd0}, 1'h0};
  assign T_3540 = T_3248 ? s2_data_2 : {{63'd0}, 1'h0};
  assign T_3542 = T_3249 ? s2_data_3 : {{63'd0}, 1'h0};
  assign T_3544 = T_3536 | T_3538;
  assign T_3545 = T_3544 | T_3540;
  assign T_3546 = T_3545 | T_3542;
  assign s2_data_muxed = T_3546;
  assign T_3553_0 = s2_data_muxed;
  assign T_3560_0 = s2_data_muxed;
  assign T_3568_0 = 1'h0;
  assign T_3570 = T_3568_0 >> 1'h0;
  assign T_3574 = s2_sc_fail == 1'h0;
  assign T_3575 = T_3445 & T_3574;
  assign T_3583 = T_3575 & T_3342;
  assign amoalu_clk = clk;
  assign amoalu_reset = reset;
  assign amoalu_io_addr = s2_req_addr[5:0];
  assign amoalu_io_cmd = s2_req_cmd;
  assign amoalu_io_typ = s2_req_typ;
  assign amoalu_io_lhs = s2_data_word;
  assign amoalu_io_rhs = s2_req_data;
  assign T_3584 = s2_valid | s2_replay;
  assign T_3592 = T_3342 | T_3570;
  assign T_3593 = T_3584 & T_3592;
  assign T_3594 = T_3570 ? T_3553_0 : amoalu_io_out;
  assign GEN_51 = T_3593 ? s2_req_addr : s3_req_addr;
  assign GEN_52 = T_3593 ? s2_req_tag : s3_req_tag;
  assign GEN_53 = T_3593 ? s2_req_cmd : s3_req_cmd;
  assign GEN_54 = T_3593 ? s2_req_typ : s3_req_typ;
  assign GEN_55 = T_3593 ? s2_req_phys : s3_req_phys;
  assign GEN_56 = T_3593 ? T_3594 : s3_req_data;
  assign GEN_57 = T_3593 ? s2_tag_match_way : s3_way;
  assign GEN_92 = {{1'd0}, 1'h1};
  assign rowWMask = GEN_92 << 1'h0;
  assign T_3598 = T_5872;
  assign T_3602 = T_3601[0];
  assign T_3603 = T_3601[2];
  assign T_3604 = T_3602 ^ T_3603;
  assign T_3605 = T_3601[3];
  assign T_3606 = T_3604 ^ T_3605;
  assign T_3607 = T_3601[5];
  assign T_3608 = T_3606 ^ T_3607;
  assign T_3609 = T_3601[15:1];
  assign T_3610 = {T_3608,T_3609};
  assign GEN_58 = T_3598 ? T_3610 : T_3601;
  assign T_3611 = T_3601[1:0];
  assign s1_replaced_way_en = GEN_85 << T_3611;
  assign GEN_59 = s1_clk_en ? T_3611 : T_3614;
  assign s2_replaced_way_en = GEN_85 << T_3614;
  assign T_3616 = s1_replaced_way_en[0];
  assign T_3617 = s1_clk_en & T_3616;
  assign GEN_60 = T_3617 ? meta_io_resp_0_tag : T_3618_tag;
  assign GEN_61 = T_3617 ? meta_io_resp_0_coh_state : T_3618_coh_state;
  assign T_3714 = s1_replaced_way_en[1];
  assign T_3715 = s1_clk_en & T_3714;
  assign GEN_62 = T_3715 ? meta_io_resp_1_tag : T_3716_tag;
  assign GEN_63 = T_3715 ? meta_io_resp_1_coh_state : T_3716_coh_state;
  assign T_3812 = s1_replaced_way_en[2];
  assign T_3813 = s1_clk_en & T_3812;
  assign GEN_64 = T_3813 ? meta_io_resp_2_tag : T_3814_tag;
  assign GEN_65 = T_3813 ? meta_io_resp_2_coh_state : T_3814_coh_state;
  assign T_3910 = s1_replaced_way_en[3];
  assign T_3911 = s1_clk_en & T_3910;
  assign GEN_66 = T_3911 ? meta_io_resp_3_tag : T_3912_tag;
  assign GEN_67 = T_3911 ? meta_io_resp_3_coh_state : T_3912_coh_state;
  assign T_4773_0_tag = T_3618_tag;
  assign T_4773_0_coh_state = T_3618_coh_state;
  assign T_4773_1_tag = T_3716_tag;
  assign T_4773_1_coh_state = T_3716_coh_state;
  assign T_4773_2_tag = T_3814_tag;
  assign T_4773_2_coh_state = T_3814_coh_state;
  assign T_4773_3_tag = T_3912_tag;
  assign T_4773_3_coh_state = T_3912_coh_state;
  assign T_5250 = s2_replaced_way_en[0];
  assign T_5251 = s2_replaced_way_en[1];
  assign T_5252 = s2_replaced_way_en[2];
  assign T_5253 = s2_replaced_way_en[3];
  assign T_5254 = {T_4773_0_tag,T_4773_0_coh_state};
  assign T_5256 = T_5250 ? T_5254 : {{21'd0}, 1'h0};
  assign T_5257 = {T_4773_1_tag,T_4773_1_coh_state};
  assign T_5259 = T_5251 ? T_5257 : {{21'd0}, 1'h0};
  assign T_5260 = {T_4773_2_tag,T_4773_2_coh_state};
  assign T_5262 = T_5252 ? T_5260 : {{21'd0}, 1'h0};
  assign T_5263 = {T_4773_3_tag,T_4773_3_coh_state};
  assign T_5265 = T_5253 ? T_5263 : {{21'd0}, 1'h0};
  assign T_5362 = T_5256 | T_5259;
  assign T_5363 = T_5362 | T_5262;
  assign T_5364 = T_5363 | T_5265;
  assign s2_repl_meta_tag = T_5557;
  assign s2_repl_meta_coh_state = T_5556;
  assign T_5556 = T_5364[1:0];
  assign T_5557 = T_5364[21:2];
  assign T_5559 = s2_hit == 1'h0;
  assign T_5560 = s2_valid_masked & T_5559;
  assign T_5561 = s2_req_cmd == 5'h2;
  assign T_5563 = T_5561 | T_3343;
  assign T_5564 = s2_req_cmd == 5'h0;
  assign T_5566 = T_5564 | T_3345;
  assign T_5568 = T_5566 | T_3337;
  assign T_5572 = T_5568 | T_3341;
  assign T_5573 = T_5563 | T_5572;
  assign T_5581 = T_5573 | T_3342;
  assign T_5582 = T_5560 & T_5581;
  assign T_5679_tag = s2_repl_meta_tag;
  assign T_5679_coh_state = s2_hit_state_state;
  assign T_5775_tag = s2_tag_match ? T_5679_tag : s2_repl_meta_tag;
  assign T_5775_coh_state = s2_tag_match ? T_5679_coh_state : s2_repl_meta_coh_state;
  assign T_5871 = s2_tag_match ? s2_tag_match_way : s2_replaced_way_en;
  assign T_5872 = mshrs_io_req_ready & mshrs_io_req_valid;
  assign T_5876 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign releaseArb_clk = clk;
  assign releaseArb_reset = reset;
  assign releaseArb_io_in_0_valid = wb_io_release_valid;
  assign releaseArb_io_in_0_bits_addr_beat = wb_io_release_bits_addr_beat;
  assign releaseArb_io_in_0_bits_addr_block = wb_io_release_bits_addr_block;
  assign releaseArb_io_in_0_bits_client_xact_id = wb_io_release_bits_client_xact_id;
  assign releaseArb_io_in_0_bits_voluntary = wb_io_release_bits_voluntary;
  assign releaseArb_io_in_0_bits_r_type = wb_io_release_bits_r_type;
  assign releaseArb_io_in_0_bits_data = wb_io_release_bits_data;
  assign releaseArb_io_in_1_valid = prober_io_rep_valid;
  assign releaseArb_io_in_1_bits_addr_beat = prober_io_rep_bits_addr_beat;
  assign releaseArb_io_in_1_bits_addr_block = prober_io_rep_bits_addr_block;
  assign releaseArb_io_in_1_bits_client_xact_id = prober_io_rep_bits_client_xact_id;
  assign releaseArb_io_in_1_bits_voluntary = prober_io_rep_bits_voluntary;
  assign releaseArb_io_in_1_bits_r_type = prober_io_rep_bits_r_type;
  assign releaseArb_io_in_1_bits_data = prober_io_rep_bits_data;
  assign releaseArb_io_out_ready = io_mem_release_ready;
  assign T_5909 = io_mem_probe_valid & T_3447;
  assign T_5912 = prober_io_req_ready & T_3447;
  assign FlowThroughSerializer_1_1_clk = clk;
  assign FlowThroughSerializer_1_1_reset = reset;
  assign FlowThroughSerializer_1_1_io_in_valid = io_mem_grant_valid;
  assign FlowThroughSerializer_1_1_io_in_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign FlowThroughSerializer_1_1_io_in_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign FlowThroughSerializer_1_1_io_in_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign FlowThroughSerializer_1_1_io_in_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign FlowThroughSerializer_1_1_io_in_bits_g_type = io_mem_grant_bits_g_type;
  assign FlowThroughSerializer_1_1_io_in_bits_data = io_mem_grant_bits_data;
  assign FlowThroughSerializer_1_1_io_in_bits_manager_id = io_mem_grant_bits_manager_id;
  assign FlowThroughSerializer_1_1_io_out_ready = T_5943;
  assign T_5913 = FlowThroughSerializer_1_1_io_out_ready & FlowThroughSerializer_1_1_io_out_valid;
  assign T_5921_0 = 3'h5;
  assign T_5921_1 = 3'h4;
  assign GEN_95 = {{1'd0}, T_5921_0};
  assign T_5923 = GEN_95 == FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign GEN_96 = {{1'd0}, T_5921_1};
  assign T_5924 = GEN_96 == FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign T_5927 = T_5923 | T_5924;
  assign T_5933_0 = 2'h0;
  assign T_5933_1 = 2'h1;
  assign GEN_97 = {{2'd0}, T_5933_0};
  assign T_5935 = GEN_97 == FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign GEN_98 = {{2'd0}, T_5933_1};
  assign T_5936 = GEN_98 == FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign T_5939 = T_5935 | T_5936;
  assign T_5940 = FlowThroughSerializer_1_1_io_out_bits_is_builtin_type ? T_5927 : T_5939;
  assign T_5942 = T_5940 == 1'h0;
  assign T_5943 = writeArb_io_in_1_ready | T_5942;
  assign T_5951_0 = 3'h5;
  assign T_5951_1 = 3'h4;
  assign GEN_99 = {{1'd0}, T_5951_0};
  assign T_5953 = GEN_99 == FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign GEN_100 = {{1'd0}, T_5951_1};
  assign T_5954 = GEN_100 == FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign T_5957 = T_5953 | T_5954;
  assign T_5963_0 = 2'h0;
  assign T_5963_1 = 2'h1;
  assign GEN_101 = {{2'd0}, T_5963_0};
  assign T_5965 = GEN_101 == FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign GEN_102 = {{2'd0}, T_5963_1};
  assign T_5966 = GEN_102 == FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign T_5969 = T_5965 | T_5966;
  assign T_5970 = FlowThroughSerializer_1_1_io_out_bits_is_builtin_type ? T_5957 : T_5969;
  assign T_5971 = FlowThroughSerializer_1_1_io_out_valid & T_5970;
  assign T_5973 = FlowThroughSerializer_1_1_io_out_bits_client_xact_id < 2'h2;
  assign T_5974 = T_5971 & T_5973;
  assign T_5977 = FlowThroughSerializer_1_1_io_out_bits_data;
  assign T_5979 = FlowThroughSerializer_1_1_io_out_valid == 1'h0;
  assign T_5980 = T_5979 | FlowThroughSerializer_1_1_io_out_ready;
  assign wbArb_clk = clk;
  assign wbArb_reset = reset;
  assign wbArb_io_in_0_valid = prober_io_wb_req_valid;
  assign wbArb_io_in_0_bits_addr_beat = prober_io_wb_req_bits_addr_beat;
  assign wbArb_io_in_0_bits_addr_block = prober_io_wb_req_bits_addr_block;
  assign wbArb_io_in_0_bits_client_xact_id = prober_io_wb_req_bits_client_xact_id;
  assign wbArb_io_in_0_bits_voluntary = prober_io_wb_req_bits_voluntary;
  assign wbArb_io_in_0_bits_r_type = prober_io_wb_req_bits_r_type;
  assign wbArb_io_in_0_bits_data = prober_io_wb_req_bits_data;
  assign wbArb_io_in_0_bits_way_en = prober_io_wb_req_bits_way_en;
  assign wbArb_io_in_1_valid = mshrs_io_wb_req_valid;
  assign wbArb_io_in_1_bits_addr_beat = mshrs_io_wb_req_bits_addr_beat;
  assign wbArb_io_in_1_bits_addr_block = mshrs_io_wb_req_bits_addr_block;
  assign wbArb_io_in_1_bits_client_xact_id = mshrs_io_wb_req_bits_client_xact_id;
  assign wbArb_io_in_1_bits_voluntary = mshrs_io_wb_req_bits_voluntary;
  assign wbArb_io_in_1_bits_r_type = mshrs_io_wb_req_bits_r_type;
  assign wbArb_io_in_1_bits_data = mshrs_io_wb_req_bits_data;
  assign wbArb_io_in_1_bits_way_en = mshrs_io_wb_req_bits_way_en;
  assign wbArb_io_out_ready = wb_io_req_ready;
  assign T_6036 = s3_valid & metaReadArb_io_out_valid;
  assign GEN_69 = T_6036 ? s3_req_addr : s4_req_addr;
  assign GEN_70 = T_6036 ? s3_req_tag : s4_req_tag;
  assign GEN_71 = T_6036 ? s3_req_cmd : s4_req_cmd;
  assign GEN_72 = T_6036 ? s3_req_typ : s4_req_typ;
  assign GEN_73 = T_6036 ? s3_req_phys : s4_req_phys;
  assign GEN_74 = T_6036 ? s3_req_data : s4_req_data;
  assign T_6112 = s2_valid_masked | s2_replay;
  assign T_6115 = T_6112 & T_3574;
  assign T_6116 = s1_addr[31:3];
  assign T_6117 = s2_req_addr[39:3];
  assign GEN_103 = {{8'd0}, T_6116};
  assign T_6118 = GEN_103 == T_6117;
  assign T_6119 = T_6115 & T_6118;
  assign T_6127 = T_6119 & T_3342;
  assign T_6129 = s3_req_addr[39:3];
  assign T_6130 = GEN_103 == T_6129;
  assign T_6131 = s3_valid & T_6130;
  assign T_6132 = s3_req_cmd == 5'h1;
  assign T_6133 = s3_req_cmd == 5'h7;
  assign T_6134 = T_6132 | T_6133;
  assign T_6135 = s3_req_cmd[3];
  assign T_6136 = s3_req_cmd == 5'h4;
  assign T_6137 = T_6135 | T_6136;
  assign T_6138 = T_6134 | T_6137;
  assign T_6139 = T_6131 & T_6138;
  assign T_6141 = s4_req_addr[39:3];
  assign T_6142 = GEN_103 == T_6141;
  assign T_6143 = s4_valid & T_6142;
  assign T_6144 = s4_req_cmd == 5'h1;
  assign T_6145 = s4_req_cmd == 5'h7;
  assign T_6146 = T_6144 | T_6145;
  assign T_6147 = s4_req_cmd[3];
  assign T_6148 = s4_req_cmd == 5'h4;
  assign T_6149 = T_6147 | T_6148;
  assign T_6150 = T_6146 | T_6149;
  assign T_6151 = T_6143 & T_6150;
  assign T_6155 = T_6127 | T_6139;
  assign T_6156 = T_6155 | T_6151;
  assign T_6157 = T_6139 ? s3_req_data : s4_req_data;
  assign T_6158 = T_6127 ? amoalu_io_out : T_6157;
  assign GEN_75 = T_6156 ? T_6158 : s2_store_bypass_data;
  assign GEN_77 = s1_clk_en ? T_6156 : s2_store_bypass;
  assign GEN_78 = s1_clk_en ? GEN_75 : s2_store_bypass_data;
  assign s2_data_word_prebypass = T_3560_0 >> 7'h0;
  assign s2_data_word = s2_store_bypass ? s2_store_bypass_data : s2_data_word_prebypass;
  assign T_6162 = s2_req_typ[1:0];
  assign T_6163 = $signed(s2_req_typ);
  assign GEN_106 = $signed(1'h0);
  assign GEN_107 = {3{GEN_106}};
  assign T_6165 = $signed(T_6163) >= $signed(GEN_107);
  assign T_6166 = dtlb_io_req_valid & dtlb_io_resp_miss;
  assign T_6167 = s1_req_addr[11:6];
  assign T_6168 = T_6167 == prober_io_meta_write_bits_idx;
  assign T_6170 = prober_io_req_ready == 1'h0;
  assign T_6171 = T_6168 & T_6170;
  assign s1_nack = T_6166 | T_6171;
  assign T_6172 = s1_valid | s1_replay;
  assign GEN_79 = T_6172 ? s1_nack : s2_nack_hit;
  assign GEN_80 = s2_nack_hit ? 1'h0 : T_5582;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T_6177 = mshrs_io_req_ready == 1'h0;
  assign s2_nack_miss = T_5559 & T_6177;
  assign T_6178 = s2_nack_hit | s2_nack_victim;
  assign s2_nack = T_6178 | s2_nack_miss;
  assign T_6180 = s2_nack == 1'h0;
  assign T_6181 = s2_valid & T_6180;
  assign T_6183 = T_3584 & s2_hit;
  assign s2_recycle_ecc = T_6183 & T_3570;
  assign GEN_81 = T_6172 ? s2_recycle_ecc : s2_recycle_next;
  assign T_6186 = s2_recycle_ecc | s2_recycle_next;
  assign T_6188 = s2_valid | block_miss;
  assign T_6189 = T_6188 & s2_nack_miss;
  assign GEN_82 = block_miss ? 1'h0 : GEN_33;
  assign cache_resp_valid = T_6593;
  assign cache_resp_bits_addr = s2_req_addr;
  assign cache_resp_bits_tag = s2_req_tag;
  assign cache_resp_bits_cmd = s2_req_cmd;
  assign cache_resp_bits_typ = s2_req_typ;
  assign cache_resp_bits_data = T_6660;
  assign cache_resp_bits_replay = s2_replay;
  assign cache_resp_bits_has_data = T_5572;
  assign cache_resp_bits_data_word_bypass = GEN_93;
  assign cache_resp_bits_store_data = s2_req_data;
  assign T_6590 = s2_replay | T_3444;
  assign T_6592 = T_3570 == 1'h0;
  assign T_6593 = T_6590 & T_6592;
  assign T_6603 = s2_req_addr[2];
  assign T_6604 = s2_data_word[63:32];
  assign T_6605 = s2_data_word[31:0];
  assign T_6606 = T_6603 ? T_6604 : T_6605;
  assign T_6612 = T_6162 == 2'h2;
  assign T_6614 = T_6606[31];
  assign T_6615 = T_6165 & T_6614;
  assign GEN_108 = {{31'd0}, T_6615};
  assign T_6617 = 32'h0 - GEN_108;
  assign T_6618 = T_6617[31:0];
  assign T_6620 = T_6612 ? T_6618 : T_6604;
  assign T_6621 = {T_6620,T_6606};
  assign T_6622 = s2_req_addr[1];
  assign T_6623 = T_6621[31:16];
  assign T_6624 = T_6621[15:0];
  assign T_6625 = T_6622 ? T_6623 : T_6624;
  assign T_6631 = T_6162 == GEN_92;
  assign T_6633 = T_6625[15];
  assign T_6634 = T_6165 & T_6633;
  assign GEN_110 = {{47'd0}, T_6634};
  assign T_6636 = 48'h0 - GEN_110;
  assign T_6637 = T_6636[47:0];
  assign T_6638 = T_6621[63:16];
  assign T_6639 = T_6631 ? T_6637 : T_6638;
  assign T_6640 = {T_6639,T_6625};
  assign T_6641 = s2_req_addr[0];
  assign T_6642 = T_6640[15:8];
  assign T_6643 = T_6640[7:0];
  assign T_6644 = T_6641 ? T_6642 : T_6643;
  assign T_6648 = T_3337 ? {{7'd0}, 1'h0} : T_6644;
  assign GEN_111 = {{1'd0}, 1'h0};
  assign T_6650 = T_6162 == GEN_111;
  assign T_6651 = T_6650 | T_3337;
  assign T_6652 = T_6648[7];
  assign T_6653 = T_6165 & T_6652;
  assign GEN_112 = {{55'd0}, T_6653};
  assign T_6655 = 56'h0 - GEN_112;
  assign T_6656 = T_6655[55:0];
  assign T_6657 = T_6640[63:8];
  assign T_6658 = T_6651 ? T_6656 : T_6657;
  assign T_6659 = {T_6658,T_6648};
  assign GEN_113 = {{63'd0}, s2_sc_fail};
  assign T_6660 = T_6659 | GEN_113;
  assign uncache_resp_valid = mshrs_io_resp_valid;
  assign uncache_resp_bits_addr = mshrs_io_resp_bits_addr;
  assign uncache_resp_bits_tag = mshrs_io_resp_bits_tag;
  assign uncache_resp_bits_cmd = mshrs_io_resp_bits_cmd;
  assign uncache_resp_bits_typ = mshrs_io_resp_bits_typ;
  assign uncache_resp_bits_data = mshrs_io_resp_bits_data;
  assign uncache_resp_bits_replay = mshrs_io_resp_bits_replay;
  assign uncache_resp_bits_has_data = mshrs_io_resp_bits_has_data;
  assign uncache_resp_bits_data_word_bypass = mshrs_io_resp_bits_data_word_bypass;
  assign uncache_resp_bits_store_data = mshrs_io_resp_bits_store_data;
  assign T_7061 = T_6172 == 1'h0;
  assign T_7063 = s2_valid & s2_nack;
  assign T_7064_valid = mshrs_io_resp_ready ? uncache_resp_valid : cache_resp_valid;
  assign T_7064_bits_addr = mshrs_io_resp_ready ? uncache_resp_bits_addr : cache_resp_bits_addr;
  assign T_7064_bits_tag = mshrs_io_resp_ready ? uncache_resp_bits_tag : cache_resp_bits_tag;
  assign T_7064_bits_cmd = mshrs_io_resp_ready ? uncache_resp_bits_cmd : cache_resp_bits_cmd;
  assign T_7064_bits_typ = mshrs_io_resp_ready ? uncache_resp_bits_typ : cache_resp_bits_typ;
  assign T_7064_bits_data = mshrs_io_resp_ready ? uncache_resp_bits_data : cache_resp_bits_data;
  assign T_7064_bits_replay = mshrs_io_resp_ready ? uncache_resp_bits_replay : cache_resp_bits_replay;
  assign T_7064_bits_has_data = mshrs_io_resp_ready ? uncache_resp_bits_has_data : cache_resp_bits_has_data;
  assign T_7064_bits_store_data = mshrs_io_resp_ready ? uncache_resp_bits_store_data : cache_resp_bits_store_data;
  assign T_7245 = mshrs_io_fence_rdy & T_2822;
  assign T_7247 = s2_valid == 1'h0;
  assign T_7248 = T_7245 & T_7247;
  assign T_7249 = s1_replay & s1_read;
  assign T_7250 = T_7249 | mshrs_io_replay_next;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_94 = {1{$random}};
  s1_valid = GEN_94[0:0];
  GEN_104 = {2{$random}};
  s1_req_addr = GEN_104[39:0];
  GEN_105 = {1{$random}};
  s1_req_tag = GEN_105[8:0];
  GEN_109 = {1{$random}};
  s1_req_cmd = GEN_109[4:0];
  GEN_114 = {1{$random}};
  s1_req_typ = GEN_114[2:0];
  GEN_115 = {1{$random}};
  s1_req_phys = GEN_115[0:0];
  GEN_116 = {2{$random}};
  s1_req_data = GEN_116[63:0];
  GEN_117 = {1{$random}};
  s1_replay = GEN_117[0:0];
  GEN_118 = {1{$random}};
  s1_clk_en = GEN_118[0:0];
  GEN_119 = {1{$random}};
  s2_valid = GEN_119[0:0];
  GEN_120 = {2{$random}};
  s2_req_addr = GEN_120[39:0];
  GEN_121 = {1{$random}};
  s2_req_tag = GEN_121[8:0];
  GEN_122 = {1{$random}};
  s2_req_cmd = GEN_122[4:0];
  GEN_123 = {1{$random}};
  s2_req_typ = GEN_123[2:0];
  GEN_124 = {1{$random}};
  s2_req_phys = GEN_124[0:0];
  GEN_125 = {2{$random}};
  s2_req_data = GEN_125[63:0];
  GEN_126 = {1{$random}};
  T_2239 = GEN_126[0:0];
  GEN_127 = {1{$random}};
  s3_valid = GEN_127[0:0];
  GEN_128 = {2{$random}};
  s3_req_addr = GEN_128[39:0];
  GEN_129 = {1{$random}};
  s3_req_tag = GEN_129[8:0];
  GEN_130 = {1{$random}};
  s3_req_cmd = GEN_130[4:0];
  GEN_131 = {1{$random}};
  s3_req_typ = GEN_131[2:0];
  GEN_132 = {1{$random}};
  s3_req_phys = GEN_132[0:0];
  GEN_133 = {2{$random}};
  s3_req_data = GEN_133[63:0];
  GEN_134 = {1{$random}};
  s3_way = GEN_134[3:0];
  GEN_135 = {1{$random}};
  s1_recycled = GEN_135[0:0];
  GEN_136 = {1{$random}};
  T_2373 = GEN_136[0:0];
  GEN_137 = {1{$random}};
  s2_tag_match_way = GEN_137[3:0];
  GEN_138 = {1{$random}};
  T_2827_state = GEN_138[1:0];
  GEN_139 = {1{$random}};
  T_2852_state = GEN_139[1:0];
  GEN_140 = {1{$random}};
  T_2877_state = GEN_140[1:0];
  GEN_141 = {1{$random}};
  T_2902_state = GEN_141[1:0];
  GEN_142 = {1{$random}};
  lrsc_count = GEN_142[4:0];
  GEN_143 = {2{$random}};
  lrsc_addr = GEN_143[33:0];
  GEN_144 = {2{$random}};
  T_3465_0 = GEN_144[63:0];
  GEN_145 = {2{$random}};
  T_3483_0 = GEN_145[63:0];
  GEN_146 = {2{$random}};
  T_3501_0 = GEN_146[63:0];
  GEN_147 = {2{$random}};
  T_3519_0 = GEN_147[63:0];
  GEN_148 = {1{$random}};
  T_3601 = GEN_148[15:0];
  GEN_149 = {1{$random}};
  T_3614 = GEN_149[1:0];
  GEN_150 = {1{$random}};
  T_3618_tag = GEN_150[19:0];
  GEN_151 = {1{$random}};
  T_3618_coh_state = GEN_151[1:0];
  GEN_152 = {1{$random}};
  T_3716_tag = GEN_152[19:0];
  GEN_153 = {1{$random}};
  T_3716_coh_state = GEN_153[1:0];
  GEN_154 = {1{$random}};
  T_3814_tag = GEN_154[19:0];
  GEN_155 = {1{$random}};
  T_3814_coh_state = GEN_155[1:0];
  GEN_156 = {1{$random}};
  T_3912_tag = GEN_156[19:0];
  GEN_157 = {1{$random}};
  T_3912_coh_state = GEN_157[1:0];
  GEN_158 = {1{$random}};
  s4_valid = GEN_158[0:0];
  GEN_159 = {2{$random}};
  s4_req_addr = GEN_159[39:0];
  GEN_160 = {1{$random}};
  s4_req_tag = GEN_160[8:0];
  GEN_161 = {1{$random}};
  s4_req_cmd = GEN_161[4:0];
  GEN_162 = {1{$random}};
  s4_req_typ = GEN_162[2:0];
  GEN_163 = {1{$random}};
  s4_req_phys = GEN_163[0:0];
  GEN_164 = {2{$random}};
  s4_req_data = GEN_164[63:0];
  GEN_165 = {2{$random}};
  s2_store_bypass_data = GEN_165[63:0];
  GEN_166 = {1{$random}};
  s2_store_bypass = GEN_166[0:0];
  GEN_167 = {1{$random}};
  s2_nack_hit = GEN_167[0:0];
  GEN_168 = {1{$random}};
  s2_recycle_next = GEN_168[0:0];
  GEN_169 = {1{$random}};
  block_miss = GEN_169[0:0];
  GEN_170 = {1{$random}};
  T_7062 = GEN_170[0:0];
  GEN_171 = {1{$random}};
  GEN_68 = GEN_171[1:0];
  GEN_172 = {1{$random}};
  GEN_76 = GEN_172[3:0];
  GEN_173 = {1{$random}};
  GEN_86 = GEN_173[3:0];
  GEN_174 = {2{$random}};
  GEN_93 = GEN_174[63:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_2081;
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_addr <= s2_req_addr;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_addr <= mshrs_io_replay_bits_addr;
        end else begin
          if(prober_io_meta_read_valid) begin
            s1_req_addr <= {{8'd0}, T_2352};
          end else begin
            if(wb_io_meta_read_valid) begin
              s1_req_addr <= {{8'd0}, T_2349};
            end else begin
              if(io_cpu_req_valid) begin
                s1_req_addr <= io_cpu_req_bits_addr;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_tag <= s2_req_tag;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_tag <= mshrs_io_replay_bits_tag;
        end else begin
          if(io_cpu_req_valid) begin
            s1_req_tag <= io_cpu_req_bits_tag;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_cmd <= s2_req_cmd;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_cmd <= mshrs_io_replay_bits_cmd;
        end else begin
          if(io_cpu_req_valid) begin
            s1_req_cmd <= io_cpu_req_bits_cmd;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_typ <= s2_req_typ;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_typ <= mshrs_io_replay_bits_typ;
        end else begin
          if(io_cpu_req_valid) begin
            s1_req_typ <= io_cpu_req_bits_typ;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_phys <= s2_req_phys;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_phys <= mshrs_io_replay_bits_phys;
        end else begin
          if(prober_io_meta_read_valid) begin
            s1_req_phys <= 1'h1;
          end else begin
            if(wb_io_meta_read_valid) begin
              s1_req_phys <= 1'h1;
            end else begin
              if(io_cpu_req_valid) begin
                s1_req_phys <= io_cpu_req_bits_phys;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_data <= s2_req_data;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_data <= mshrs_io_replay_bits_data;
        end else begin
          if(io_cpu_req_valid) begin
            s1_req_data <= io_cpu_req_bits_data;
          end
        end
      end
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T_5876;
    end
    if(1'h0) begin
    end else begin
      s1_clk_en <= metaReadArb_io_out_valid;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_addr <= {{8'd0}, s1_addr};
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_tag <= s1_req_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_typ <= s1_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_phys <= s1_req_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        if(s1_recycled) begin
          s2_req_data <= s1_req_data;
        end else begin
          if(s1_write) begin
            if(s1_replay) begin
              s2_req_data <= mshrs_io_replay_bits_data;
            end else begin
              s2_req_data <= io_cpu_s1_data;
            end
          end
        end
      end
    end
    if(reset) begin
      T_2239 <= 1'h0;
    end else begin
      T_2239 <= s1_replay;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T_3583;
    end
    if(1'h0) begin
    end else begin
      if(T_3593) begin
        s3_req_addr <= s2_req_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3593) begin
        s3_req_tag <= s2_req_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3593) begin
        s3_req_cmd <= s2_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3593) begin
        s3_req_typ <= s2_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3593) begin
        s3_req_phys <= s2_req_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3593) begin
        if(T_3570) begin
          s3_req_data <= T_3553_0;
        end else begin
          s3_req_data <= amoalu_io_out;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3593) begin
        s3_way <= s2_tag_match_way;
      end
    end
    if(reset) begin
      s1_recycled <= 1'h0;
    end else begin
      if(s1_clk_en) begin
        s1_recycled <= s2_recycle;
      end
    end
    if(1'h0) begin
    end else begin
      T_2373 <= T_2372;
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_tag_match_way <= s1_tag_match_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_2827_state <= meta_io_resp_0_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_2852_state <= meta_io_resp_1_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_2877_state <= meta_io_resp_2_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_2902_state <= meta_io_resp_3_coh_state;
      end
    end
    if(reset) begin
      lrsc_count <= {{4'd0}, 1'h0};
    end else begin
      if(io_cpu_invalidate_lr) begin
        lrsc_count <= {{4'd0}, 1'h0};
      end else begin
        if(T_3445) begin
          if(T_3337) begin
            lrsc_count <= {{4'd0}, 1'h0};
          end else begin
            if(T_3345) begin
              if(T_3447) begin
                lrsc_count <= 5'h1f;
              end else begin
                if(lrsc_valid) begin
                  lrsc_count <= T_3443;
                end
              end
            end else begin
              if(lrsc_valid) begin
                lrsc_count <= T_3443;
              end
            end
          end
        end else begin
          if(lrsc_valid) begin
            lrsc_count <= T_3443;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3445) begin
        if(T_3345) begin
          lrsc_addr <= T_2780;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3468) begin
        T_3465_0 <= T_3476;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3486) begin
        T_3483_0 <= T_3494;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3504) begin
        T_3501_0 <= T_3512;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3522) begin
        T_3519_0 <= T_3530;
      end
    end
    if(reset) begin
      T_3601 <= 16'h1;
    end else begin
      if(T_3598) begin
        T_3601 <= T_3610;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_3614 <= T_3611;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3617) begin
        T_3618_tag <= meta_io_resp_0_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3617) begin
        T_3618_coh_state <= meta_io_resp_0_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3715) begin
        T_3716_tag <= meta_io_resp_1_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3715) begin
        T_3716_coh_state <= meta_io_resp_1_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3813) begin
        T_3814_tag <= meta_io_resp_2_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3813) begin
        T_3814_coh_state <= meta_io_resp_2_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3911) begin
        T_3912_tag <= meta_io_resp_3_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3911) begin
        T_3912_coh_state <= meta_io_resp_3_coh_state;
      end
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(1'h0) begin
    end else begin
      if(T_6036) begin
        s4_req_addr <= s3_req_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_6036) begin
        s4_req_tag <= s3_req_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_6036) begin
        s4_req_cmd <= s3_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_6036) begin
        s4_req_typ <= s3_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_6036) begin
        s4_req_phys <= s3_req_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_6036) begin
        s4_req_data <= s3_req_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        if(T_6156) begin
          if(T_6127) begin
            s2_store_bypass_data <= amoalu_io_out;
          end else begin
            if(T_6139) begin
              s2_store_bypass_data <= s3_req_data;
            end else begin
              s2_store_bypass_data <= s4_req_data;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_store_bypass <= T_6156;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_6172) begin
        s2_nack_hit <= s1_nack;
      end
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else begin
      if(T_6172) begin
        s2_recycle_next <= s2_recycle_ecc;
      end
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T_6189;
    end
    if(1'h0) begin
    end else begin
      T_7062 <= T_7061;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2379) begin
          $fwrite(32'h80000002,"Assertion failed: DCache exception occurred - cache response not killed.\n    at nbdcache.scala:866 assert (!(Reg(next=\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2379) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_2379) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOArbiter(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output [2:0] io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [1:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [1:0] io_out_grant_bits_client_xact_id,
  input  [2:0] io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module RRArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [26:0] io_in_0_bits_addr,
  input  [1:0] io_in_0_bits_prv,
  input   io_in_0_bits_store,
  input   io_in_0_bits_fetch,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [26:0] io_in_1_bits_addr,
  input  [1:0] io_in_1_bits_prv,
  input   io_in_1_bits_store,
  input   io_in_1_bits_fetch,
  input   io_out_ready,
  output  io_out_valid,
  output [26:0] io_out_bits_addr,
  output [1:0] io_out_bits_prv,
  output  io_out_bits_store,
  output  io_out_bits_fetch,
  output  io_chosen
);
  wire  T_143;
  wire  GEN_0;
  wire  GEN_5;
  wire [26:0] GEN_1;
  wire [26:0] GEN_6;
  wire [1:0] GEN_2;
  wire [1:0] GEN_7;
  wire  GEN_3;
  wire  GEN_8;
  wire  GEN_4;
  wire  GEN_9;
  wire  T_169;
  reg  T_170;
  reg [31:0] GEN_13;
  wire  GEN_10;
  wire  T_173;
  wire  T_175;
  wire  T_178;
  wire  T_182;
  wire  T_184;
  wire  T_188;
  wire  T_189;
  wire  T_190;
  wire  GEN_11;
  wire  GEN_12;
  assign io_in_0_ready = T_189;
  assign io_in_1_ready = T_190;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr = GEN_1;
  assign io_out_bits_prv = GEN_2;
  assign io_out_bits_store = GEN_3;
  assign io_out_bits_fetch = GEN_4;
  assign io_chosen = T_143;
  assign T_143 = GEN_12;
  assign GEN_0 = GEN_5;
  assign GEN_5 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_6;
  assign GEN_6 = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign GEN_2 = GEN_7;
  assign GEN_7 = io_chosen ? io_in_1_bits_prv : io_in_0_bits_prv;
  assign GEN_3 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_bits_store : io_in_0_bits_store;
  assign GEN_4 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_fetch : io_in_0_bits_fetch;
  assign T_169 = io_out_ready & io_out_valid;
  assign GEN_10 = T_169 ? io_chosen : T_170;
  assign T_173 = 1'h1 > T_170;
  assign T_175 = io_in_1_valid & T_173;
  assign T_178 = T_175 | io_in_0_valid;
  assign T_182 = T_175 == 1'h0;
  assign T_184 = T_178 == 1'h0;
  assign T_188 = T_173 | T_184;
  assign T_189 = T_182 & io_out_ready;
  assign T_190 = T_188 & io_out_ready;
  assign GEN_11 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_12 = T_175 ? 1'h1 : GEN_11;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_13 = {1{$random}};
  T_170 = GEN_13[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_169) begin
        T_170 <= io_chosen;
      end
    end
  end
endmodule
module PTW(
  input   clk,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [26:0] io_requestor_0_req_bits_addr,
  input  [1:0] io_requestor_0_req_bits_prv,
  input   io_requestor_0_req_bits_store,
  input   io_requestor_0_req_bits_fetch,
  output  io_requestor_0_resp_valid,
  output [19:0] io_requestor_0_resp_bits_pte_ppn,
  output [2:0] io_requestor_0_resp_bits_pte_reserved_for_software,
  output  io_requestor_0_resp_bits_pte_d,
  output  io_requestor_0_resp_bits_pte_r,
  output [3:0] io_requestor_0_resp_bits_pte_typ,
  output  io_requestor_0_resp_bits_pte_v,
  output [6:0] io_requestor_0_ptbr_asid,
  output [37:0] io_requestor_0_ptbr_ppn,
  output  io_requestor_0_invalidate,
  output  io_requestor_0_status_debug,
  output [1:0] io_requestor_0_status_prv,
  output  io_requestor_0_status_sd,
  output [30:0] io_requestor_0_status_zero3,
  output  io_requestor_0_status_sd_rv32,
  output [1:0] io_requestor_0_status_zero2,
  output [4:0] io_requestor_0_status_vm,
  output [4:0] io_requestor_0_status_zero1,
  output  io_requestor_0_status_pum,
  output  io_requestor_0_status_mprv,
  output [1:0] io_requestor_0_status_xs,
  output [1:0] io_requestor_0_status_fs,
  output [1:0] io_requestor_0_status_mpp,
  output [1:0] io_requestor_0_status_hpp,
  output  io_requestor_0_status_spp,
  output  io_requestor_0_status_mpie,
  output  io_requestor_0_status_hpie,
  output  io_requestor_0_status_spie,
  output  io_requestor_0_status_upie,
  output  io_requestor_0_status_mie,
  output  io_requestor_0_status_hie,
  output  io_requestor_0_status_sie,
  output  io_requestor_0_status_uie,
  output  io_requestor_1_req_ready,
  input   io_requestor_1_req_valid,
  input  [26:0] io_requestor_1_req_bits_addr,
  input  [1:0] io_requestor_1_req_bits_prv,
  input   io_requestor_1_req_bits_store,
  input   io_requestor_1_req_bits_fetch,
  output  io_requestor_1_resp_valid,
  output [19:0] io_requestor_1_resp_bits_pte_ppn,
  output [2:0] io_requestor_1_resp_bits_pte_reserved_for_software,
  output  io_requestor_1_resp_bits_pte_d,
  output  io_requestor_1_resp_bits_pte_r,
  output [3:0] io_requestor_1_resp_bits_pte_typ,
  output  io_requestor_1_resp_bits_pte_v,
  output [6:0] io_requestor_1_ptbr_asid,
  output [37:0] io_requestor_1_ptbr_ppn,
  output  io_requestor_1_invalidate,
  output  io_requestor_1_status_debug,
  output [1:0] io_requestor_1_status_prv,
  output  io_requestor_1_status_sd,
  output [30:0] io_requestor_1_status_zero3,
  output  io_requestor_1_status_sd_rv32,
  output [1:0] io_requestor_1_status_zero2,
  output [4:0] io_requestor_1_status_vm,
  output [4:0] io_requestor_1_status_zero1,
  output  io_requestor_1_status_pum,
  output  io_requestor_1_status_mprv,
  output [1:0] io_requestor_1_status_xs,
  output [1:0] io_requestor_1_status_fs,
  output [1:0] io_requestor_1_status_mpp,
  output [1:0] io_requestor_1_status_hpp,
  output  io_requestor_1_status_spp,
  output  io_requestor_1_status_mpie,
  output  io_requestor_1_status_hpie,
  output  io_requestor_1_status_spie,
  output  io_requestor_1_status_upie,
  output  io_requestor_1_status_mie,
  output  io_requestor_1_status_hie,
  output  io_requestor_1_status_sie,
  output  io_requestor_1_status_uie,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [8:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [63:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [63:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,
  input  [39:0] io_mem_resp_bits_addr,
  input  [8:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,
  input  [63:0] io_mem_resp_bits_data,
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input  [63:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered,
  input  [6:0] io_dpath_ptbr_asid,
  input  [37:0] io_dpath_ptbr_ppn,
  input   io_dpath_invalidate,
  input   io_dpath_status_debug,
  input  [1:0] io_dpath_status_prv,
  input   io_dpath_status_sd,
  input  [30:0] io_dpath_status_zero3,
  input   io_dpath_status_sd_rv32,
  input  [1:0] io_dpath_status_zero2,
  input  [4:0] io_dpath_status_vm,
  input  [4:0] io_dpath_status_zero1,
  input   io_dpath_status_pum,
  input   io_dpath_status_mprv,
  input  [1:0] io_dpath_status_xs,
  input  [1:0] io_dpath_status_fs,
  input  [1:0] io_dpath_status_mpp,
  input  [1:0] io_dpath_status_hpp,
  input   io_dpath_status_spp,
  input   io_dpath_status_mpie,
  input   io_dpath_status_hpie,
  input   io_dpath_status_spie,
  input   io_dpath_status_upie,
  input   io_dpath_status_mie,
  input   io_dpath_status_hie,
  input   io_dpath_status_sie,
  input   io_dpath_status_uie
);
  reg [2:0] state;
  reg [31:0] GEN_20;
  reg [1:0] count;
  reg [31:0] GEN_21;
  reg [26:0] r_req_addr;
  reg [31:0] GEN_22;
  reg [1:0] r_req_prv;
  reg [31:0] GEN_23;
  reg  r_req_store;
  reg [31:0] GEN_24;
  reg  r_req_fetch;
  reg [31:0] GEN_25;
  reg  r_req_dest;
  reg [31:0] GEN_26;
  reg [19:0] r_pte_ppn;
  reg [31:0] GEN_27;
  reg [2:0] r_pte_reserved_for_software;
  reg [31:0] GEN_28;
  reg  r_pte_d;
  reg [31:0] GEN_41;
  reg  r_pte_r;
  reg [31:0] GEN_42;
  reg [3:0] r_pte_typ;
  reg [31:0] GEN_73;
  reg  r_pte_v;
  reg [31:0] GEN_75;
  wire [8:0] T_1910;
  wire [17:0] T_1912;
  wire [8:0] T_1913;
  wire [8:0] T_1915;
  wire [8:0] T_1921_0;
  wire [8:0] T_1921_1;
  wire [8:0] T_1921_2;
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [26:0] arb_io_in_0_bits_addr;
  wire [1:0] arb_io_in_0_bits_prv;
  wire  arb_io_in_0_bits_store;
  wire  arb_io_in_0_bits_fetch;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [26:0] arb_io_in_1_bits_addr;
  wire [1:0] arb_io_in_1_bits_prv;
  wire  arb_io_in_1_bits_store;
  wire  arb_io_in_1_bits_fetch;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [26:0] arb_io_out_bits_addr;
  wire [1:0] arb_io_out_bits_prv;
  wire  arb_io_out_bits_store;
  wire  arb_io_out_bits_fetch;
  wire  arb_io_chosen;
  wire  T_1928;
  wire [19:0] pte_ppn;
  wire [2:0] pte_reserved_for_software;
  wire  pte_d;
  wire  pte_r;
  wire [3:0] pte_typ;
  wire  pte_v;
  wire  T_1949;
  wire [3:0] T_1950;
  wire  T_1951;
  wire  T_1952;
  wire [2:0] T_1953;
  wire [19:0] T_1954;
  wire [8:0] GEN_0;
  wire [1:0] GEN_69;
  wire [8:0] GEN_4;
  wire [8:0] GEN_5;
  wire [28:0] T_1955;
  wire [31:0] GEN_70;
  wire [31:0] pte_addr;
  wire  T_1956;
  wire [26:0] GEN_6;
  wire [1:0] GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [37:0] GEN_11;
  reg [2:0] T_1958;
  reg [31:0] GEN_80;
  reg  T_1965_0;
  reg [31:0] GEN_81;
  reg  T_1965_1;
  reg [31:0] GEN_82;
  reg  T_1965_2;
  reg [31:0] GEN_83;
  wire [1:0] T_1967;
  wire [2:0] T_1968;
  reg [31:0] T_1971 [0:2];
  reg [31:0] GEN_84;
  wire [31:0] T_1971_T_1976_data;
  wire [1:0] T_1971_T_1976_addr;
  wire  T_1971_T_1976_en;
  wire [31:0] T_1971_T_1979_data;
  wire [1:0] T_1971_T_1979_addr;
  wire  T_1971_T_1979_en;
  wire [31:0] T_1971_T_1982_data;
  wire [1:0] T_1971_T_1982_addr;
  wire  T_1971_T_1982_en;
  wire [31:0] T_1971_T_2024_data;
  wire [1:0] T_1971_T_2024_addr;
  wire  T_1971_T_2024_mask;
  wire  T_1971_T_2024_en;
  reg [19:0] T_1974 [0:2];
  reg [31:0] GEN_85;
  wire [19:0] T_1974_T_2064_data;
  wire [1:0] T_1974_T_2064_addr;
  wire  T_1974_T_2064_en;
  wire [19:0] T_1974_T_2066_data;
  wire [1:0] T_1974_T_2066_addr;
  wire  T_1974_T_2066_en;
  wire [19:0] T_1974_T_2068_data;
  wire [1:0] T_1974_T_2068_addr;
  wire  T_1974_T_2068_en;
  wire [19:0] T_1974_T_2025_data;
  wire [1:0] T_1974_T_2025_addr;
  wire  T_1974_T_2025_mask;
  wire  T_1974_T_2025_en;
  wire  T_1977;
  wire  T_1980;
  wire  T_1983;
  wire  T_1989_0;
  wire  T_1989_1;
  wire  T_1989_2;
  wire [1:0] T_1991;
  wire [2:0] T_1992;
  wire [2:0] T_1993;
  wire [2:0] GEN_71;
  wire  pte_cache_hit;
  wire [3:0] GEN_72;
  wire  T_1996;
  wire  T_1997;
  wire  T_1998;
  wire  T_2000;
  wire  T_2001;
  wire [2:0] T_2002;
  wire  T_2004;
  wire [2:0] T_2006;
  wire  T_2007;
  wire [1:0] T_2008;
  wire [2:0] T_2009;
  wire  T_2010;
  wire [2:0] T_2011;
  wire [1:0] T_2012;
  wire  T_2014;
  wire  T_2015;
  wire [1:0] T_2020;
  wire [1:0] T_2021;
  wire [1:0] T_2022;
  wire  GEN_1;
  wire [1:0] GEN_74;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  T_2026;
  wire  T_2027;
  wire  T_2028;
  wire [1:0] T_2029;
  wire [1:0] GEN_76;
  wire [1:0] T_2032;
  wire  T_2033;
  wire [1:0] T_2034;
  wire  T_2036;
  wire [3:0] GEN_77;
  wire [3:0] T_2038;
  wire [2:0] T_2039;
  wire [2:0] T_2040;
  wire [2:0] T_2041;
  wire [2:0] T_2043;
  wire [2:0] T_2044;
  wire [1:0] T_2045;
  wire  T_2046;
  wire [5:0] GEN_78;
  wire [5:0] T_2048;
  wire [2:0] T_2049;
  wire [2:0] T_2050;
  wire [2:0] T_2051;
  wire [2:0] T_2053;
  wire [2:0] T_2054;
  wire [2:0] GEN_29;
  wire  T_2056;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  T_2060;
  wire  T_2061;
  wire [19:0] T_2070;
  wire [19:0] T_2072;
  wire [19:0] T_2074;
  wire [19:0] T_2076;
  wire [19:0] T_2077;
  wire [19:0] pte_cache_data;
  wire  T_2078;
  wire [3:0] GEN_79;
  wire  T_2080;
  wire  T_2081;
  wire  T_2082;
  wire  T_2083;
  wire  T_2085;
  wire  T_2086;
  wire  T_2087;
  wire  T_2088;
  wire  T_2092;
  wire  T_2093;
  wire  T_2098;
  wire  T_2099;
  wire  T_2101;
  wire  T_2109;
  wire  T_2116;
  wire  T_2117;
  wire  perm_ok;
  wire  T_2119;
  wire  T_2121;
  wire  T_2122;
  wire  T_2123;
  wire  set_dirty_bit;
  wire  T_2124;
  wire  T_2125;
  wire  T_2127;
  wire  T_2128;
  wire [37:0] GEN_33;
  wire [2:0] GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [3:0] GEN_37;
  wire  GEN_38;
  wire [19:0] T_2144_ppn;
  wire [2:0] T_2144_reserved_for_software;
  wire  T_2144_d;
  wire  T_2144_r;
  wire [3:0] T_2144_typ;
  wire  T_2144_v;
  wire [29:0] T_2152;
  wire  T_2153;
  wire [3:0] T_2154;
  wire  T_2155;
  wire  T_2156;
  wire [2:0] T_2157;
  wire [19:0] T_2158;
  wire [19:0] pte_wdata_ppn;
  wire [2:0] pte_wdata_reserved_for_software;
  wire  pte_wdata_d;
  wire  pte_wdata_r;
  wire [3:0] pte_wdata_typ;
  wire  pte_wdata_v;
  wire  T_2167;
  wire  T_2168;
  wire [4:0] T_2171;
  wire [4:0] T_2172;
  wire [5:0] T_2173;
  wire [22:0] T_2174;
  wire [23:0] T_2175;
  wire [29:0] T_2176;
  wire [27:0] r_resp_ppn;
  wire [9:0] T_2179;
  wire [17:0] T_2180;
  wire [27:0] T_2181;
  wire [18:0] T_2182;
  wire [27:0] T_2184;
  wire [27:0] T_2190_0;
  wire [27:0] T_2190_1;
  wire [27:0] T_2190_2;
  wire  resp_val;
  wire  T_2193;
  wire  T_2194;
  wire [27:0] GEN_2;
  wire [27:0] GEN_39;
  wire [27:0] GEN_40;
  wire  T_2197;
  wire [27:0] GEN_3;
  wire  T_2198;
  wire [2:0] GEN_43;
  wire [2:0] GEN_44;
  wire [1:0] GEN_45;
  wire  T_2200;
  wire  T_2202;
  wire  T_2203;
  wire [2:0] T_2206;
  wire [1:0] T_2207;
  wire  GEN_46;
  wire [2:0] GEN_47;
  wire [1:0] GEN_48;
  wire [37:0] GEN_49;
  wire  T_2209;
  wire  T_2210;
  wire [2:0] GEN_50;
  wire  GEN_51;
  wire [2:0] GEN_52;
  wire [1:0] GEN_53;
  wire [37:0] GEN_54;
  wire  T_2211;
  wire [2:0] GEN_55;
  wire  T_2215;
  wire [2:0] GEN_56;
  wire  T_2221;
  wire [2:0] GEN_57;
  wire [1:0] GEN_58;
  wire [2:0] GEN_59;
  wire [1:0] GEN_60;
  wire [2:0] GEN_61;
  wire [1:0] GEN_62;
  wire  T_2225;
  wire [2:0] GEN_63;
  wire [2:0] GEN_64;
  wire  T_2226;
  wire [2:0] GEN_65;
  wire [2:0] GEN_66;
  wire [2:0] GEN_67;
  wire  T_2227;
  wire [2:0] GEN_68;
  reg [8:0] GEN_15;
  reg [31:0] GEN_86;
  reg [63:0] GEN_19;
  reg [63:0] GEN_87;
  RRArbiter arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_prv(arb_io_in_0_bits_prv),
    .io_in_0_bits_store(arb_io_in_0_bits_store),
    .io_in_0_bits_fetch(arb_io_in_0_bits_fetch),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_prv(arb_io_in_1_bits_prv),
    .io_in_1_bits_store(arb_io_in_1_bits_store),
    .io_in_1_bits_fetch(arb_io_in_1_bits_fetch),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_prv(arb_io_out_bits_prv),
    .io_out_bits_store(arb_io_out_bits_store),
    .io_out_bits_fetch(arb_io_out_bits_fetch),
    .io_chosen(arb_io_chosen)
  );
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_0_resp_valid = T_2194;
  assign io_requestor_0_resp_bits_pte_ppn = GEN_2[19:0];
  assign io_requestor_0_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_0_resp_bits_pte_d = r_pte_d;
  assign io_requestor_0_resp_bits_pte_r = r_pte_r;
  assign io_requestor_0_resp_bits_pte_typ = r_pte_typ;
  assign io_requestor_0_resp_bits_pte_v = r_pte_v;
  assign io_requestor_0_ptbr_asid = io_dpath_ptbr_asid;
  assign io_requestor_0_ptbr_ppn = io_dpath_ptbr_ppn;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_debug = io_dpath_status_debug;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_sd = io_dpath_status_sd;
  assign io_requestor_0_status_zero3 = io_dpath_status_zero3;
  assign io_requestor_0_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_0_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_0_status_pum = io_dpath_status_pum;
  assign io_requestor_0_status_mprv = io_dpath_status_mprv;
  assign io_requestor_0_status_xs = io_dpath_status_xs;
  assign io_requestor_0_status_fs = io_dpath_status_fs;
  assign io_requestor_0_status_mpp = io_dpath_status_mpp;
  assign io_requestor_0_status_hpp = io_dpath_status_hpp;
  assign io_requestor_0_status_spp = io_dpath_status_spp;
  assign io_requestor_0_status_mpie = io_dpath_status_mpie;
  assign io_requestor_0_status_hpie = io_dpath_status_hpie;
  assign io_requestor_0_status_spie = io_dpath_status_spie;
  assign io_requestor_0_status_upie = io_dpath_status_upie;
  assign io_requestor_0_status_mie = io_dpath_status_mie;
  assign io_requestor_0_status_hie = io_dpath_status_hie;
  assign io_requestor_0_status_sie = io_dpath_status_sie;
  assign io_requestor_0_status_uie = io_dpath_status_uie;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  assign io_requestor_1_resp_valid = T_2197;
  assign io_requestor_1_resp_bits_pte_ppn = GEN_3[19:0];
  assign io_requestor_1_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_1_resp_bits_pte_d = r_pte_d;
  assign io_requestor_1_resp_bits_pte_r = r_pte_r;
  assign io_requestor_1_resp_bits_pte_typ = r_pte_typ;
  assign io_requestor_1_resp_bits_pte_v = r_pte_v;
  assign io_requestor_1_ptbr_asid = io_dpath_ptbr_asid;
  assign io_requestor_1_ptbr_ppn = io_dpath_ptbr_ppn;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_debug = io_dpath_status_debug;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_sd = io_dpath_status_sd;
  assign io_requestor_1_status_zero3 = io_dpath_status_zero3;
  assign io_requestor_1_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_1_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_1_status_pum = io_dpath_status_pum;
  assign io_requestor_1_status_mprv = io_dpath_status_mprv;
  assign io_requestor_1_status_xs = io_dpath_status_xs;
  assign io_requestor_1_status_fs = io_dpath_status_fs;
  assign io_requestor_1_status_mpp = io_dpath_status_mpp;
  assign io_requestor_1_status_hpp = io_dpath_status_hpp;
  assign io_requestor_1_status_spp = io_dpath_status_spp;
  assign io_requestor_1_status_mpie = io_dpath_status_mpie;
  assign io_requestor_1_status_hpie = io_dpath_status_hpie;
  assign io_requestor_1_status_spie = io_dpath_status_spie;
  assign io_requestor_1_status_upie = io_dpath_status_upie;
  assign io_requestor_1_status_mie = io_dpath_status_mie;
  assign io_requestor_1_status_hie = io_dpath_status_hie;
  assign io_requestor_1_status_sie = io_dpath_status_sie;
  assign io_requestor_1_status_uie = io_dpath_status_uie;
  assign io_mem_req_valid = GEN_51;
  assign io_mem_req_bits_addr = {{8'd0}, pte_addr};
  assign io_mem_req_bits_tag = GEN_15;
  assign io_mem_req_bits_cmd = T_2171;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_data = GEN_19;
  assign io_mem_s1_kill = 1'h0;
  assign io_mem_s1_data = {{34'd0}, T_2176};
  assign io_mem_invalidate_lr = 1'h0;
  assign T_1910 = r_req_addr[26:18];
  assign T_1912 = r_req_addr[26:9];
  assign T_1913 = T_1912[8:0];
  assign T_1915 = r_req_addr[8:0];
  assign T_1921_0 = T_1910;
  assign T_1921_1 = T_1913;
  assign T_1921_2 = T_1915;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_requestor_0_req_valid;
  assign arb_io_in_0_bits_addr = io_requestor_0_req_bits_addr;
  assign arb_io_in_0_bits_prv = io_requestor_0_req_bits_prv;
  assign arb_io_in_0_bits_store = io_requestor_0_req_bits_store;
  assign arb_io_in_0_bits_fetch = io_requestor_0_req_bits_fetch;
  assign arb_io_in_1_valid = io_requestor_1_req_valid;
  assign arb_io_in_1_bits_addr = io_requestor_1_req_bits_addr;
  assign arb_io_in_1_bits_prv = io_requestor_1_req_bits_prv;
  assign arb_io_in_1_bits_store = io_requestor_1_req_bits_store;
  assign arb_io_in_1_bits_fetch = io_requestor_1_req_bits_fetch;
  assign arb_io_out_ready = T_1928;
  assign T_1928 = state == 3'h0;
  assign pte_ppn = T_1954;
  assign pte_reserved_for_software = T_1953;
  assign pte_d = T_1952;
  assign pte_r = T_1951;
  assign pte_typ = T_1950;
  assign pte_v = T_1949;
  assign T_1949 = io_mem_resp_bits_data[0];
  assign T_1950 = io_mem_resp_bits_data[4:1];
  assign T_1951 = io_mem_resp_bits_data[5];
  assign T_1952 = io_mem_resp_bits_data[6];
  assign T_1953 = io_mem_resp_bits_data[9:7];
  assign T_1954 = io_mem_resp_bits_data[29:10];
  assign GEN_0 = GEN_5;
  assign GEN_69 = {{1'd0}, 1'h1};
  assign GEN_4 = GEN_69 == count ? T_1921_1 : T_1921_0;
  assign GEN_5 = 2'h2 == count ? T_1921_2 : GEN_4;
  assign T_1955 = {r_pte_ppn,GEN_0};
  assign GEN_70 = {{3'd0}, T_1955};
  assign pte_addr = GEN_70 << 3;
  assign T_1956 = arb_io_out_ready & arb_io_out_valid;
  assign GEN_6 = T_1956 ? arb_io_out_bits_addr : r_req_addr;
  assign GEN_7 = T_1956 ? arb_io_out_bits_prv : r_req_prv;
  assign GEN_8 = T_1956 ? arb_io_out_bits_store : r_req_store;
  assign GEN_9 = T_1956 ? arb_io_out_bits_fetch : r_req_fetch;
  assign GEN_10 = T_1956 ? arb_io_chosen : r_req_dest;
  assign GEN_11 = T_1956 ? io_dpath_ptbr_ppn : {{18'd0}, r_pte_ppn};
  assign T_1967 = {T_1965_2,T_1965_1};
  assign T_1968 = {T_1967,T_1965_0};
  assign T_1971_T_1976_addr = {{1'd0}, 1'h0};
  assign T_1971_T_1976_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1971_T_1976_data = T_1971[T_1971_T_1976_addr];
  `else
  assign T_1971_T_1976_data = T_1971_T_1976_addr >= 2'h3 ? $random : T_1971[T_1971_T_1976_addr];
  `endif
  assign T_1971_T_1979_addr = {{1'd0}, 1'h1};
  assign T_1971_T_1979_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1971_T_1979_data = T_1971[T_1971_T_1979_addr];
  `else
  assign T_1971_T_1979_data = T_1971_T_1979_addr >= 2'h3 ? $random : T_1971[T_1971_T_1979_addr];
  `endif
  assign T_1971_T_1982_addr = 2'h2;
  assign T_1971_T_1982_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1971_T_1982_data = T_1971[T_1971_T_1982_addr];
  `else
  assign T_1971_T_1982_data = T_1971_T_1982_addr >= 2'h3 ? $random : T_1971[T_1971_T_1982_addr];
  `endif
  assign T_1971_T_2024_data = pte_addr;
  assign T_1971_T_2024_addr = T_2022;
  assign T_1971_T_2024_mask = T_2001;
  assign T_1971_T_2024_en = T_2001;
  assign T_1974_T_2064_addr = {{1'd0}, 1'h0};
  assign T_1974_T_2064_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1974_T_2064_data = T_1974[T_1974_T_2064_addr];
  `else
  assign T_1974_T_2064_data = T_1974_T_2064_addr >= 2'h3 ? $random : T_1974[T_1974_T_2064_addr];
  `endif
  assign T_1974_T_2066_addr = {{1'd0}, 1'h1};
  assign T_1974_T_2066_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1974_T_2066_data = T_1974[T_1974_T_2066_addr];
  `else
  assign T_1974_T_2066_data = T_1974_T_2066_addr >= 2'h3 ? $random : T_1974[T_1974_T_2066_addr];
  `endif
  assign T_1974_T_2068_addr = 2'h2;
  assign T_1974_T_2068_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1974_T_2068_data = T_1974[T_1974_T_2068_addr];
  `else
  assign T_1974_T_2068_data = T_1974_T_2068_addr >= 2'h3 ? $random : T_1974[T_1974_T_2068_addr];
  `endif
  assign T_1974_T_2025_data = pte_ppn;
  assign T_1974_T_2025_addr = T_2022;
  assign T_1974_T_2025_mask = T_2001;
  assign T_1974_T_2025_en = T_2001;
  assign T_1977 = T_1971_T_1976_data == pte_addr;
  assign T_1980 = T_1971_T_1979_data == pte_addr;
  assign T_1983 = T_1971_T_1982_data == pte_addr;
  assign T_1989_0 = T_1977;
  assign T_1989_1 = T_1980;
  assign T_1989_2 = T_1983;
  assign T_1991 = {T_1989_2,T_1989_1};
  assign T_1992 = {T_1991,T_1989_0};
  assign T_1993 = T_1992 & T_1968;
  assign GEN_71 = {{2'd0}, 1'h0};
  assign pte_cache_hit = T_1993 != GEN_71;
  assign GEN_72 = {{2'd0}, 2'h2};
  assign T_1996 = pte_typ < GEN_72;
  assign T_1997 = pte_v & T_1996;
  assign T_1998 = io_mem_resp_valid & T_1997;
  assign T_2000 = pte_cache_hit == 1'h0;
  assign T_2001 = T_1998 & T_2000;
  assign T_2002 = ~ T_1968;
  assign T_2004 = T_2002 == GEN_71;
  assign T_2006 = T_1958 >> 1'h1;
  assign T_2007 = T_2006[0];
  assign T_2008 = {1'h1,T_2007};
  assign T_2009 = T_1958 >> T_2008;
  assign T_2010 = T_2009[0];
  assign T_2011 = {T_2008,T_2010};
  assign T_2012 = T_2011[1:0];
  assign T_2014 = T_2002[0];
  assign T_2015 = T_2002[1];
  assign T_2020 = T_2015 ? {{1'd0}, 1'h1} : 2'h2;
  assign T_2021 = T_2014 ? {{1'd0}, 1'h0} : T_2020;
  assign T_2022 = T_2004 ? T_2012 : T_2021;
  assign GEN_1 = 1'h1;
  assign GEN_74 = {{1'd0}, 1'h0};
  assign GEN_12 = GEN_74 == T_2022 ? GEN_1 : T_1965_0;
  assign GEN_13 = GEN_69 == T_2022 ? GEN_1 : T_1965_1;
  assign GEN_14 = 2'h2 == T_2022 ? GEN_1 : T_1965_2;
  assign GEN_16 = T_2001 ? GEN_12 : T_1965_0;
  assign GEN_17 = T_2001 ? GEN_13 : T_1965_1;
  assign GEN_18 = T_2001 ? GEN_14 : T_1965_2;
  assign T_2026 = state == 3'h1;
  assign T_2027 = pte_cache_hit & T_2026;
  assign T_2028 = T_1993[2];
  assign T_2029 = T_1993[1:0];
  assign GEN_76 = {{1'd0}, T_2028};
  assign T_2032 = GEN_76 | T_2029;
  assign T_2033 = T_2032[1];
  assign T_2034 = {T_2028,T_2033};
  assign T_2036 = T_2034[1];
  assign GEN_77 = {{1'd0}, 3'h1};
  assign T_2038 = GEN_77 << 1'h1;
  assign T_2039 = T_2038[2:0];
  assign T_2040 = ~ T_2039;
  assign T_2041 = T_1958 & T_2040;
  assign T_2043 = T_2036 ? {{2'd0}, 1'h0} : T_2039;
  assign T_2044 = T_2041 | T_2043;
  assign T_2045 = {1'h1,T_2036};
  assign T_2046 = T_2034[0];
  assign GEN_78 = {{3'd0}, 3'h1};
  assign T_2048 = GEN_78 << T_2045;
  assign T_2049 = T_2048[2:0];
  assign T_2050 = ~ T_2049;
  assign T_2051 = T_2044 & T_2050;
  assign T_2053 = T_2046 ? {{2'd0}, 1'h0} : T_2049;
  assign T_2054 = T_2051 | T_2053;
  assign GEN_29 = T_2027 ? T_2054 : T_1958;
  assign T_2056 = reset | io_dpath_invalidate;
  assign GEN_30 = T_2056 ? 1'h0 : GEN_16;
  assign GEN_31 = T_2056 ? 1'h0 : GEN_17;
  assign GEN_32 = T_2056 ? 1'h0 : GEN_18;
  assign T_2060 = T_1993[0];
  assign T_2061 = T_1993[1];
  assign T_2070 = T_2060 ? T_1974_T_2064_data : {{19'd0}, 1'h0};
  assign T_2072 = T_2061 ? T_1974_T_2066_data : {{19'd0}, 1'h0};
  assign T_2074 = T_2028 ? T_1974_T_2068_data : {{19'd0}, 1'h0};
  assign T_2076 = T_2070 | T_2072;
  assign T_2077 = T_2076 | T_2074;
  assign pte_cache_data = T_2077;
  assign T_2078 = r_req_prv[0];
  assign GEN_79 = {{1'd0}, 3'h4};
  assign T_2080 = pte_typ >= GEN_79;
  assign T_2081 = pte_v & T_2080;
  assign T_2082 = pte_typ[1];
  assign T_2083 = T_2081 & T_2082;
  assign T_2085 = pte_typ >= GEN_72;
  assign T_2086 = pte_v & T_2085;
  assign T_2087 = pte_typ[0];
  assign T_2088 = T_2086 & T_2087;
  assign T_2092 = r_req_store ? T_2088 : T_2086;
  assign T_2093 = r_req_fetch ? T_2083 : T_2092;
  assign T_2098 = pte_typ < 4'h8;
  assign T_2099 = T_2086 & T_2098;
  assign T_2101 = T_2099 & T_2082;
  assign T_2109 = T_2099 & T_2087;
  assign T_2116 = r_req_store ? T_2109 : T_2099;
  assign T_2117 = r_req_fetch ? T_2101 : T_2116;
  assign perm_ok = T_2078 ? T_2093 : T_2117;
  assign T_2119 = pte_r == 1'h0;
  assign T_2121 = pte_d == 1'h0;
  assign T_2122 = r_req_store & T_2121;
  assign T_2123 = T_2119 | T_2122;
  assign set_dirty_bit = perm_ok & T_2123;
  assign T_2124 = state == 3'h2;
  assign T_2125 = io_mem_resp_valid & T_2124;
  assign T_2127 = set_dirty_bit == 1'h0;
  assign T_2128 = T_2125 & T_2127;
  assign GEN_33 = T_2128 ? {{18'd0}, pte_ppn} : GEN_11;
  assign GEN_34 = T_2128 ? pte_reserved_for_software : r_pte_reserved_for_software;
  assign GEN_35 = T_2128 ? pte_d : r_pte_d;
  assign GEN_36 = T_2128 ? pte_r : r_pte_r;
  assign GEN_37 = T_2128 ? pte_typ : r_pte_typ;
  assign GEN_38 = T_2128 ? pte_v : r_pte_v;
  assign T_2144_ppn = T_2158;
  assign T_2144_reserved_for_software = T_2157;
  assign T_2144_d = T_2156;
  assign T_2144_r = T_2155;
  assign T_2144_typ = T_2154;
  assign T_2144_v = T_2153;
  assign T_2152 = {{29'd0}, 1'h0};
  assign T_2153 = T_2152[0];
  assign T_2154 = T_2152[4:1];
  assign T_2155 = T_2152[5];
  assign T_2156 = T_2152[6];
  assign T_2157 = T_2152[9:7];
  assign T_2158 = T_2152[29:10];
  assign pte_wdata_ppn = T_2144_ppn;
  assign pte_wdata_reserved_for_software = T_2144_reserved_for_software;
  assign pte_wdata_d = r_req_store;
  assign pte_wdata_r = 1'h1;
  assign pte_wdata_typ = T_2144_typ;
  assign pte_wdata_v = T_2144_v;
  assign T_2167 = state == 3'h3;
  assign T_2168 = T_2026 | T_2167;
  assign T_2171 = T_2167 ? 5'ha : 5'h0;
  assign T_2172 = {pte_wdata_r,pte_wdata_typ};
  assign T_2173 = {T_2172,pte_wdata_v};
  assign T_2174 = {pte_wdata_ppn,pte_wdata_reserved_for_software};
  assign T_2175 = {T_2174,pte_wdata_d};
  assign T_2176 = {T_2175,T_2173};
  assign r_resp_ppn = io_mem_req_bits_addr[39:12];
  assign T_2179 = r_resp_ppn[27:18];
  assign T_2180 = r_req_addr[17:0];
  assign T_2181 = {T_2179,T_2180};
  assign T_2182 = r_resp_ppn[27:9];
  assign T_2184 = {T_2182,T_1915};
  assign T_2190_0 = T_2181;
  assign T_2190_1 = T_2184;
  assign T_2190_2 = r_resp_ppn;
  assign resp_val = state == 3'h5;
  assign T_2193 = r_req_dest == 1'h0;
  assign T_2194 = resp_val & T_2193;
  assign GEN_2 = GEN_40;
  assign GEN_39 = GEN_69 == count ? T_2190_1 : T_2190_0;
  assign GEN_40 = 2'h2 == count ? T_2190_2 : GEN_39;
  assign T_2197 = resp_val & r_req_dest;
  assign GEN_3 = GEN_40;
  assign T_2198 = 3'h0 == state;
  assign GEN_43 = arb_io_out_valid ? 3'h1 : state;
  assign GEN_44 = T_2198 ? GEN_43 : state;
  assign GEN_45 = T_2198 ? {{1'd0}, 1'h0} : count;
  assign T_2200 = 3'h1 == state;
  assign T_2202 = count < 2'h2;
  assign T_2203 = pte_cache_hit & T_2202;
  assign T_2206 = count + GEN_69;
  assign T_2207 = T_2206[1:0];
  assign GEN_46 = T_2203 ? 1'h0 : T_2168;
  assign GEN_47 = T_2203 ? 3'h1 : GEN_44;
  assign GEN_48 = T_2203 ? T_2207 : GEN_45;
  assign GEN_49 = T_2203 ? {{18'd0}, pte_cache_data} : GEN_33;
  assign T_2209 = T_2203 == 1'h0;
  assign T_2210 = T_2209 & io_mem_req_ready;
  assign GEN_50 = T_2210 ? 3'h2 : GEN_47;
  assign GEN_51 = T_2200 ? GEN_46 : T_2168;
  assign GEN_52 = T_2200 ? GEN_50 : GEN_44;
  assign GEN_53 = T_2200 ? GEN_48 : GEN_45;
  assign GEN_54 = T_2200 ? GEN_49 : GEN_33;
  assign T_2211 = 3'h2 == state;
  assign GEN_55 = io_mem_s2_nack ? 3'h1 : GEN_52;
  assign T_2215 = T_2086 & set_dirty_bit;
  assign GEN_56 = T_2215 ? 3'h3 : 3'h5;
  assign T_2221 = T_1997 & T_2202;
  assign GEN_57 = T_2221 ? 3'h1 : GEN_56;
  assign GEN_58 = T_2221 ? T_2207 : GEN_53;
  assign GEN_59 = io_mem_resp_valid ? GEN_57 : GEN_55;
  assign GEN_60 = io_mem_resp_valid ? GEN_58 : GEN_53;
  assign GEN_61 = T_2211 ? GEN_59 : GEN_52;
  assign GEN_62 = T_2211 ? GEN_60 : GEN_53;
  assign T_2225 = 3'h3 == state;
  assign GEN_63 = io_mem_req_ready ? 3'h4 : GEN_61;
  assign GEN_64 = T_2225 ? GEN_63 : GEN_61;
  assign T_2226 = 3'h4 == state;
  assign GEN_65 = io_mem_s2_nack ? 3'h3 : GEN_64;
  assign GEN_66 = io_mem_resp_valid ? 3'h1 : GEN_65;
  assign GEN_67 = T_2226 ? GEN_66 : GEN_64;
  assign T_2227 = 3'h5 == state;
  assign GEN_68 = T_2227 ? 3'h0 : GEN_67;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_20 = {1{$random}};
  state = GEN_20[2:0];
  GEN_21 = {1{$random}};
  count = GEN_21[1:0];
  GEN_22 = {1{$random}};
  r_req_addr = GEN_22[26:0];
  GEN_23 = {1{$random}};
  r_req_prv = GEN_23[1:0];
  GEN_24 = {1{$random}};
  r_req_store = GEN_24[0:0];
  GEN_25 = {1{$random}};
  r_req_fetch = GEN_25[0:0];
  GEN_26 = {1{$random}};
  r_req_dest = GEN_26[0:0];
  GEN_27 = {1{$random}};
  r_pte_ppn = GEN_27[19:0];
  GEN_28 = {1{$random}};
  r_pte_reserved_for_software = GEN_28[2:0];
  GEN_41 = {1{$random}};
  r_pte_d = GEN_41[0:0];
  GEN_42 = {1{$random}};
  r_pte_r = GEN_42[0:0];
  GEN_73 = {1{$random}};
  r_pte_typ = GEN_73[3:0];
  GEN_75 = {1{$random}};
  r_pte_v = GEN_75[0:0];
  GEN_80 = {1{$random}};
  T_1958 = GEN_80[2:0];
  GEN_81 = {1{$random}};
  T_1965_0 = GEN_81[0:0];
  GEN_82 = {1{$random}};
  T_1965_1 = GEN_82[0:0];
  GEN_83 = {1{$random}};
  T_1965_2 = GEN_83[0:0];
  GEN_84 = {1{$random}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    T_1971[initvar] = GEN_84[31:0];
  GEN_85 = {1{$random}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    T_1974[initvar] = GEN_85[19:0];
  GEN_86 = {1{$random}};
  GEN_15 = GEN_86[8:0];
  GEN_87 = {2{$random}};
  GEN_19 = GEN_87[63:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      if(T_2227) begin
        state <= 3'h0;
      end else begin
        if(T_2226) begin
          if(io_mem_resp_valid) begin
            state <= 3'h1;
          end else begin
            if(io_mem_s2_nack) begin
              state <= 3'h3;
            end else begin
              if(T_2225) begin
                if(io_mem_req_ready) begin
                  state <= 3'h4;
                end else begin
                  if(T_2211) begin
                    if(io_mem_resp_valid) begin
                      if(T_2221) begin
                        state <= 3'h1;
                      end else begin
                        if(T_2215) begin
                          state <= 3'h3;
                        end else begin
                          state <= 3'h5;
                        end
                      end
                    end else begin
                      if(io_mem_s2_nack) begin
                        state <= 3'h1;
                      end else begin
                        if(T_2200) begin
                          if(T_2210) begin
                            state <= 3'h2;
                          end else begin
                            if(T_2203) begin
                              state <= 3'h1;
                            end else begin
                              if(T_2198) begin
                                if(arb_io_out_valid) begin
                                  state <= 3'h1;
                                end
                              end
                            end
                          end
                        end else begin
                          if(T_2198) begin
                            if(arb_io_out_valid) begin
                              state <= 3'h1;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    if(T_2200) begin
                      if(T_2210) begin
                        state <= 3'h2;
                      end else begin
                        if(T_2203) begin
                          state <= 3'h1;
                        end else begin
                          if(T_2198) begin
                            if(arb_io_out_valid) begin
                              state <= 3'h1;
                            end
                          end
                        end
                      end
                    end else begin
                      if(T_2198) begin
                        if(arb_io_out_valid) begin
                          state <= 3'h1;
                        end
                      end
                    end
                  end
                end
              end else begin
                if(T_2211) begin
                  if(io_mem_resp_valid) begin
                    if(T_2221) begin
                      state <= 3'h1;
                    end else begin
                      if(T_2215) begin
                        state <= 3'h3;
                      end else begin
                        state <= 3'h5;
                      end
                    end
                  end else begin
                    if(io_mem_s2_nack) begin
                      state <= 3'h1;
                    end else begin
                      if(T_2200) begin
                        if(T_2210) begin
                          state <= 3'h2;
                        end else begin
                          if(T_2203) begin
                            state <= 3'h1;
                          end else begin
                            state <= GEN_44;
                          end
                        end
                      end else begin
                        state <= GEN_44;
                      end
                    end
                  end
                end else begin
                  if(T_2200) begin
                    if(T_2210) begin
                      state <= 3'h2;
                    end else begin
                      if(T_2203) begin
                        state <= 3'h1;
                      end else begin
                        state <= GEN_44;
                      end
                    end
                  end else begin
                    state <= GEN_44;
                  end
                end
              end
            end
          end
        end else begin
          if(T_2225) begin
            if(io_mem_req_ready) begin
              state <= 3'h4;
            end else begin
              if(T_2211) begin
                if(io_mem_resp_valid) begin
                  if(T_2221) begin
                    state <= 3'h1;
                  end else begin
                    if(T_2215) begin
                      state <= 3'h3;
                    end else begin
                      state <= 3'h5;
                    end
                  end
                end else begin
                  if(io_mem_s2_nack) begin
                    state <= 3'h1;
                  end else begin
                    state <= GEN_52;
                  end
                end
              end else begin
                state <= GEN_52;
              end
            end
          end else begin
            if(T_2211) begin
              if(io_mem_resp_valid) begin
                if(T_2221) begin
                  state <= 3'h1;
                end else begin
                  if(T_2215) begin
                    state <= 3'h3;
                  end else begin
                    state <= 3'h5;
                  end
                end
              end else begin
                if(io_mem_s2_nack) begin
                  state <= 3'h1;
                end else begin
                  state <= GEN_52;
                end
              end
            end else begin
              state <= GEN_52;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2211) begin
        if(io_mem_resp_valid) begin
          if(T_2221) begin
            count <= T_2207;
          end else begin
            if(T_2200) begin
              if(T_2203) begin
                count <= T_2207;
              end else begin
                if(T_2198) begin
                  count <= {{1'd0}, 1'h0};
                end
              end
            end else begin
              if(T_2198) begin
                count <= {{1'd0}, 1'h0};
              end
            end
          end
        end else begin
          if(T_2200) begin
            if(T_2203) begin
              count <= T_2207;
            end else begin
              if(T_2198) begin
                count <= {{1'd0}, 1'h0};
              end
            end
          end else begin
            if(T_2198) begin
              count <= {{1'd0}, 1'h0};
            end
          end
        end
      end else begin
        if(T_2200) begin
          if(T_2203) begin
            count <= T_2207;
          end else begin
            count <= GEN_45;
          end
        end else begin
          count <= GEN_45;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1956) begin
        r_req_addr <= arb_io_out_bits_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1956) begin
        r_req_prv <= arb_io_out_bits_prv;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1956) begin
        r_req_store <= arb_io_out_bits_store;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1956) begin
        r_req_fetch <= arb_io_out_bits_fetch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1956) begin
        r_req_dest <= arb_io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      r_pte_ppn <= GEN_54[19:0];
    end
    if(1'h0) begin
    end else begin
      if(T_2128) begin
        r_pte_reserved_for_software <= pte_reserved_for_software;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2128) begin
        r_pte_d <= pte_d;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2128) begin
        r_pte_r <= pte_r;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2128) begin
        r_pte_typ <= pte_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2128) begin
        r_pte_v <= pte_v;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2027) begin
        T_1958 <= T_2054;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2056) begin
        T_1965_0 <= 1'h0;
      end else begin
        if(T_2001) begin
          if(GEN_74 == T_2022) begin
            T_1965_0 <= GEN_1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2056) begin
        T_1965_1 <= 1'h0;
      end else begin
        if(T_2001) begin
          if(GEN_69 == T_2022) begin
            T_1965_1 <= GEN_1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2056) begin
        T_1965_2 <= 1'h0;
      end else begin
        if(T_2001) begin
          if(2'h2 == T_2022) begin
            T_1965_2 <= GEN_1;
          end
        end
      end
    end
    if(T_1971_T_2024_en & T_1971_T_2024_mask) begin
      T_1971[T_1971_T_2024_addr] <= T_1971_T_2024_data;
    end
    if(T_1974_T_2025_en & T_1974_T_2025_mask) begin
      T_1974[T_1974_T_2025_addr] <= T_1974_T_2025_data;
    end
  end
endmodule
module HellaCacheArbiter(
  input   clk,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [39:0] io_requestor_0_req_bits_addr,
  input  [8:0] io_requestor_0_req_bits_tag,
  input  [4:0] io_requestor_0_req_bits_cmd,
  input  [2:0] io_requestor_0_req_bits_typ,
  input   io_requestor_0_req_bits_phys,
  input  [63:0] io_requestor_0_req_bits_data,
  input   io_requestor_0_s1_kill,
  input  [63:0] io_requestor_0_s1_data,
  output  io_requestor_0_s2_nack,
  output  io_requestor_0_resp_valid,
  output [39:0] io_requestor_0_resp_bits_addr,
  output [8:0] io_requestor_0_resp_bits_tag,
  output [4:0] io_requestor_0_resp_bits_cmd,
  output [2:0] io_requestor_0_resp_bits_typ,
  output [63:0] io_requestor_0_resp_bits_data,
  output  io_requestor_0_resp_bits_replay,
  output  io_requestor_0_resp_bits_has_data,
  output [63:0] io_requestor_0_resp_bits_data_word_bypass,
  output [63:0] io_requestor_0_resp_bits_store_data,
  output  io_requestor_0_replay_next,
  output  io_requestor_0_xcpt_ma_ld,
  output  io_requestor_0_xcpt_ma_st,
  output  io_requestor_0_xcpt_pf_ld,
  output  io_requestor_0_xcpt_pf_st,
  input   io_requestor_0_invalidate_lr,
  output  io_requestor_0_ordered,
  output  io_requestor_1_req_ready,
  input   io_requestor_1_req_valid,
  input  [39:0] io_requestor_1_req_bits_addr,
  input  [8:0] io_requestor_1_req_bits_tag,
  input  [4:0] io_requestor_1_req_bits_cmd,
  input  [2:0] io_requestor_1_req_bits_typ,
  input   io_requestor_1_req_bits_phys,
  input  [63:0] io_requestor_1_req_bits_data,
  input   io_requestor_1_s1_kill,
  input  [63:0] io_requestor_1_s1_data,
  output  io_requestor_1_s2_nack,
  output  io_requestor_1_resp_valid,
  output [39:0] io_requestor_1_resp_bits_addr,
  output [8:0] io_requestor_1_resp_bits_tag,
  output [4:0] io_requestor_1_resp_bits_cmd,
  output [2:0] io_requestor_1_resp_bits_typ,
  output [63:0] io_requestor_1_resp_bits_data,
  output  io_requestor_1_resp_bits_replay,
  output  io_requestor_1_resp_bits_has_data,
  output [63:0] io_requestor_1_resp_bits_data_word_bypass,
  output [63:0] io_requestor_1_resp_bits_store_data,
  output  io_requestor_1_replay_next,
  output  io_requestor_1_xcpt_ma_ld,
  output  io_requestor_1_xcpt_ma_st,
  output  io_requestor_1_xcpt_pf_ld,
  output  io_requestor_1_xcpt_pf_st,
  input   io_requestor_1_invalidate_lr,
  output  io_requestor_1_ordered,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [8:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [63:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [63:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,
  input  [39:0] io_mem_resp_bits_addr,
  input  [8:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,
  input  [63:0] io_mem_resp_bits_data,
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input  [63:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered
);
  reg  s1_id;
  reg [31:0] GEN_9;
  reg  s2_id;
  reg [31:0] GEN_10;
  wire  T_7160;
  wire  T_7161;
  wire  T_7163;
  wire  T_7164;
  wire [9:0] T_7166;
  wire [9:0] T_7169;
  wire [4:0] GEN_0;
  wire [2:0] GEN_1;
  wire [39:0] GEN_2;
  wire  GEN_3;
  wire [9:0] GEN_4;
  wire  GEN_5;
  wire  T_7172;
  wire  GEN_6;
  wire [63:0] GEN_7;
  wire  T_7173;
  wire  T_7175;
  wire  T_7176;
  wire  T_7178;
  wire  T_7179;
  wire [7:0] T_7180;
  wire  T_7184;
  wire  T_7187;
  reg [63:0] GEN_8;
  reg [63:0] GEN_11;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_0_s2_nack = T_7179;
  assign io_requestor_0_resp_valid = T_7176;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_tag = {{1'd0}, T_7180};
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_replay_next = io_mem_replay_next;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_1_req_ready = T_7164;
  assign io_requestor_1_s2_nack = T_7187;
  assign io_requestor_1_resp_valid = T_7184;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_tag = {{1'd0}, T_7180};
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_replay_next = io_mem_replay_next;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_mem_req_valid = T_7161;
  assign io_mem_req_bits_addr = GEN_2;
  assign io_mem_req_bits_tag = GEN_4[8:0];
  assign io_mem_req_bits_cmd = GEN_0;
  assign io_mem_req_bits_typ = GEN_1;
  assign io_mem_req_bits_phys = GEN_3;
  assign io_mem_req_bits_data = GEN_8;
  assign io_mem_s1_kill = GEN_6;
  assign io_mem_s1_data = GEN_7;
  assign io_mem_invalidate_lr = T_7160;
  assign T_7160 = io_requestor_0_invalidate_lr | io_requestor_1_invalidate_lr;
  assign T_7161 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign T_7163 = io_requestor_0_req_valid == 1'h0;
  assign T_7164 = io_requestor_0_req_ready & T_7163;
  assign T_7166 = {io_requestor_1_req_bits_tag,1'h1};
  assign T_7169 = {io_requestor_0_req_bits_tag,1'h0};
  assign GEN_0 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign GEN_1 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign GEN_2 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign GEN_3 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign GEN_4 = io_requestor_0_req_valid ? T_7169 : T_7166;
  assign GEN_5 = io_requestor_0_req_valid ? 1'h0 : 1'h1;
  assign T_7172 = s1_id == 1'h0;
  assign GEN_6 = T_7172 ? io_requestor_0_s1_kill : io_requestor_1_s1_kill;
  assign GEN_7 = T_7172 ? io_requestor_0_s1_data : io_requestor_1_s1_data;
  assign T_7173 = io_mem_resp_bits_tag[0];
  assign T_7175 = T_7173 == 1'h0;
  assign T_7176 = io_mem_resp_valid & T_7175;
  assign T_7178 = s2_id == 1'h0;
  assign T_7179 = io_mem_s2_nack & T_7178;
  assign T_7180 = io_mem_resp_bits_tag[8:1];
  assign T_7184 = io_mem_resp_valid & T_7173;
  assign T_7187 = io_mem_s2_nack & s2_id;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  s1_id = GEN_9[0:0];
  GEN_10 = {1{$random}};
  s2_id = GEN_10[0:0];
  GEN_11 = {2{$random}};
  GEN_8 = GEN_11[63:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(io_requestor_0_req_valid) begin
        s1_id <= 1'h0;
      end else begin
        s1_id <= 1'h1;
      end
    end
    if(1'h0) begin
    end else begin
      s2_id <= s1_id;
    end
  end
endmodule
module RocketTile(
  input   clk,
  input   reset,
  input   io_cached_0_acquire_ready,
  output  io_cached_0_acquire_valid,
  output [25:0] io_cached_0_acquire_bits_addr_block,
  output [1:0] io_cached_0_acquire_bits_client_xact_id,
  output [2:0] io_cached_0_acquire_bits_addr_beat,
  output  io_cached_0_acquire_bits_is_builtin_type,
  output [2:0] io_cached_0_acquire_bits_a_type,
  output [11:0] io_cached_0_acquire_bits_union,
  output [63:0] io_cached_0_acquire_bits_data,
  output  io_cached_0_probe_ready,
  input   io_cached_0_probe_valid,
  input  [25:0] io_cached_0_probe_bits_addr_block,
  input  [1:0] io_cached_0_probe_bits_p_type,
  input   io_cached_0_release_ready,
  output  io_cached_0_release_valid,
  output [2:0] io_cached_0_release_bits_addr_beat,
  output [25:0] io_cached_0_release_bits_addr_block,
  output [1:0] io_cached_0_release_bits_client_xact_id,
  output  io_cached_0_release_bits_voluntary,
  output [2:0] io_cached_0_release_bits_r_type,
  output [63:0] io_cached_0_release_bits_data,
  output  io_cached_0_grant_ready,
  input   io_cached_0_grant_valid,
  input  [2:0] io_cached_0_grant_bits_addr_beat,
  input  [1:0] io_cached_0_grant_bits_client_xact_id,
  input  [2:0] io_cached_0_grant_bits_manager_xact_id,
  input   io_cached_0_grant_bits_is_builtin_type,
  input  [3:0] io_cached_0_grant_bits_g_type,
  input  [63:0] io_cached_0_grant_bits_data,
  input   io_cached_0_grant_bits_manager_id,
  input   io_cached_0_finish_ready,
  output  io_cached_0_finish_valid,
  output [2:0] io_cached_0_finish_bits_manager_xact_id,
  output  io_cached_0_finish_bits_manager_id,
  input   io_uncached_0_acquire_ready,
  output  io_uncached_0_acquire_valid,
  output [25:0] io_uncached_0_acquire_bits_addr_block,
  output [1:0] io_uncached_0_acquire_bits_client_xact_id,
  output [2:0] io_uncached_0_acquire_bits_addr_beat,
  output  io_uncached_0_acquire_bits_is_builtin_type,
  output [2:0] io_uncached_0_acquire_bits_a_type,
  output [11:0] io_uncached_0_acquire_bits_union,
  output [63:0] io_uncached_0_acquire_bits_data,
  output  io_uncached_0_grant_ready,
  input   io_uncached_0_grant_valid,
  input  [2:0] io_uncached_0_grant_bits_addr_beat,
  input  [1:0] io_uncached_0_grant_bits_client_xact_id,
  input  [2:0] io_uncached_0_grant_bits_manager_xact_id,
  input   io_uncached_0_grant_bits_is_builtin_type,
  input  [3:0] io_uncached_0_grant_bits_g_type,
  input  [63:0] io_uncached_0_grant_bits_data,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip
);
  wire  core_clk;
  wire  core_reset;
  wire  core_io_prci_reset;
  wire  core_io_prci_id;
  wire  core_io_prci_interrupts_meip;
  wire  core_io_prci_interrupts_seip;
  wire  core_io_prci_interrupts_debug;
  wire  core_io_prci_interrupts_mtip;
  wire  core_io_prci_interrupts_msip;
  wire  core_io_imem_req_valid;
  wire [39:0] core_io_imem_req_bits_pc;
  wire  core_io_imem_resp_ready;
  wire  core_io_imem_resp_valid;
  wire [39:0] core_io_imem_resp_bits_pc;
  wire [31:0] core_io_imem_resp_bits_data_0;
  wire  core_io_imem_resp_bits_mask;
  wire  core_io_imem_resp_bits_xcpt_if;
  wire  core_io_imem_btb_resp_valid;
  wire  core_io_imem_btb_resp_bits_taken;
  wire  core_io_imem_btb_resp_bits_mask;
  wire  core_io_imem_btb_resp_bits_bridx;
  wire [38:0] core_io_imem_btb_resp_bits_target;
  wire [5:0] core_io_imem_btb_resp_bits_entry;
  wire [6:0] core_io_imem_btb_resp_bits_bht_history;
  wire [1:0] core_io_imem_btb_resp_bits_bht_value;
  wire  core_io_imem_btb_update_valid;
  wire  core_io_imem_btb_update_bits_prediction_valid;
  wire  core_io_imem_btb_update_bits_prediction_bits_taken;
  wire  core_io_imem_btb_update_bits_prediction_bits_mask;
  wire  core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] core_io_imem_btb_update_bits_pc;
  wire [38:0] core_io_imem_btb_update_bits_target;
  wire  core_io_imem_btb_update_bits_taken;
  wire  core_io_imem_btb_update_bits_isJump;
  wire  core_io_imem_btb_update_bits_isReturn;
  wire [38:0] core_io_imem_btb_update_bits_br_pc;
  wire  core_io_imem_bht_update_valid;
  wire  core_io_imem_bht_update_bits_prediction_valid;
  wire  core_io_imem_bht_update_bits_prediction_bits_taken;
  wire  core_io_imem_bht_update_bits_prediction_bits_mask;
  wire  core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_bht_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] core_io_imem_bht_update_bits_pc;
  wire  core_io_imem_bht_update_bits_taken;
  wire  core_io_imem_bht_update_bits_mispredict;
  wire  core_io_imem_ras_update_valid;
  wire  core_io_imem_ras_update_bits_isCall;
  wire  core_io_imem_ras_update_bits_isReturn;
  wire [38:0] core_io_imem_ras_update_bits_returnAddr;
  wire  core_io_imem_ras_update_bits_prediction_valid;
  wire  core_io_imem_ras_update_bits_prediction_bits_taken;
  wire  core_io_imem_ras_update_bits_prediction_bits_mask;
  wire  core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_ras_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire  core_io_imem_flush_icache;
  wire  core_io_imem_flush_tlb;
  wire [39:0] core_io_imem_npc;
  wire  core_io_dmem_req_ready;
  wire  core_io_dmem_req_valid;
  wire [39:0] core_io_dmem_req_bits_addr;
  wire [8:0] core_io_dmem_req_bits_tag;
  wire [4:0] core_io_dmem_req_bits_cmd;
  wire [2:0] core_io_dmem_req_bits_typ;
  wire  core_io_dmem_req_bits_phys;
  wire [63:0] core_io_dmem_req_bits_data;
  wire  core_io_dmem_s1_kill;
  wire [63:0] core_io_dmem_s1_data;
  wire  core_io_dmem_s2_nack;
  wire  core_io_dmem_resp_valid;
  wire [39:0] core_io_dmem_resp_bits_addr;
  wire [8:0] core_io_dmem_resp_bits_tag;
  wire [4:0] core_io_dmem_resp_bits_cmd;
  wire [2:0] core_io_dmem_resp_bits_typ;
  wire [63:0] core_io_dmem_resp_bits_data;
  wire  core_io_dmem_resp_bits_replay;
  wire  core_io_dmem_resp_bits_has_data;
  wire [63:0] core_io_dmem_resp_bits_data_word_bypass;
  wire [63:0] core_io_dmem_resp_bits_store_data;
  wire  core_io_dmem_replay_next;
  wire  core_io_dmem_xcpt_ma_ld;
  wire  core_io_dmem_xcpt_ma_st;
  wire  core_io_dmem_xcpt_pf_ld;
  wire  core_io_dmem_xcpt_pf_st;
  wire  core_io_dmem_invalidate_lr;
  wire  core_io_dmem_ordered;
  wire [6:0] core_io_ptw_ptbr_asid;
  wire [37:0] core_io_ptw_ptbr_ppn;
  wire  core_io_ptw_invalidate;
  wire  core_io_ptw_status_debug;
  wire [1:0] core_io_ptw_status_prv;
  wire  core_io_ptw_status_sd;
  wire [30:0] core_io_ptw_status_zero3;
  wire  core_io_ptw_status_sd_rv32;
  wire [1:0] core_io_ptw_status_zero2;
  wire [4:0] core_io_ptw_status_vm;
  wire [4:0] core_io_ptw_status_zero1;
  wire  core_io_ptw_status_pum;
  wire  core_io_ptw_status_mprv;
  wire [1:0] core_io_ptw_status_xs;
  wire [1:0] core_io_ptw_status_fs;
  wire [1:0] core_io_ptw_status_mpp;
  wire [1:0] core_io_ptw_status_hpp;
  wire  core_io_ptw_status_spp;
  wire  core_io_ptw_status_mpie;
  wire  core_io_ptw_status_hpie;
  wire  core_io_ptw_status_spie;
  wire  core_io_ptw_status_upie;
  wire  core_io_ptw_status_mie;
  wire  core_io_ptw_status_hie;
  wire  core_io_ptw_status_sie;
  wire  core_io_ptw_status_uie;
  wire [31:0] core_io_fpu_inst;
  wire [63:0] core_io_fpu_fromint_data;
  wire [2:0] core_io_fpu_fcsr_rm;
  wire  core_io_fpu_fcsr_flags_valid;
  wire [4:0] core_io_fpu_fcsr_flags_bits;
  wire [63:0] core_io_fpu_store_data;
  wire [63:0] core_io_fpu_toint_data;
  wire  core_io_fpu_dmem_resp_val;
  wire [2:0] core_io_fpu_dmem_resp_type;
  wire [4:0] core_io_fpu_dmem_resp_tag;
  wire [63:0] core_io_fpu_dmem_resp_data;
  wire  core_io_fpu_valid;
  wire  core_io_fpu_fcsr_rdy;
  wire  core_io_fpu_nack_mem;
  wire  core_io_fpu_illegal_rm;
  wire  core_io_fpu_killx;
  wire  core_io_fpu_killm;
  wire [4:0] core_io_fpu_dec_cmd;
  wire  core_io_fpu_dec_ldst;
  wire  core_io_fpu_dec_wen;
  wire  core_io_fpu_dec_ren1;
  wire  core_io_fpu_dec_ren2;
  wire  core_io_fpu_dec_ren3;
  wire  core_io_fpu_dec_swap12;
  wire  core_io_fpu_dec_swap23;
  wire  core_io_fpu_dec_single;
  wire  core_io_fpu_dec_fromint;
  wire  core_io_fpu_dec_toint;
  wire  core_io_fpu_dec_fastpipe;
  wire  core_io_fpu_dec_fma;
  wire  core_io_fpu_dec_div;
  wire  core_io_fpu_dec_sqrt;
  wire  core_io_fpu_dec_round;
  wire  core_io_fpu_dec_wflags;
  wire  core_io_fpu_sboard_set;
  wire  core_io_fpu_sboard_clr;
  wire [4:0] core_io_fpu_sboard_clra;
  wire  core_io_fpu_cp_req_ready;
  wire  core_io_fpu_cp_req_valid;
  wire [4:0] core_io_fpu_cp_req_bits_cmd;
  wire  core_io_fpu_cp_req_bits_ldst;
  wire  core_io_fpu_cp_req_bits_wen;
  wire  core_io_fpu_cp_req_bits_ren1;
  wire  core_io_fpu_cp_req_bits_ren2;
  wire  core_io_fpu_cp_req_bits_ren3;
  wire  core_io_fpu_cp_req_bits_swap12;
  wire  core_io_fpu_cp_req_bits_swap23;
  wire  core_io_fpu_cp_req_bits_single;
  wire  core_io_fpu_cp_req_bits_fromint;
  wire  core_io_fpu_cp_req_bits_toint;
  wire  core_io_fpu_cp_req_bits_fastpipe;
  wire  core_io_fpu_cp_req_bits_fma;
  wire  core_io_fpu_cp_req_bits_div;
  wire  core_io_fpu_cp_req_bits_sqrt;
  wire  core_io_fpu_cp_req_bits_round;
  wire  core_io_fpu_cp_req_bits_wflags;
  wire [2:0] core_io_fpu_cp_req_bits_rm;
  wire [1:0] core_io_fpu_cp_req_bits_typ;
  wire [64:0] core_io_fpu_cp_req_bits_in1;
  wire [64:0] core_io_fpu_cp_req_bits_in2;
  wire [64:0] core_io_fpu_cp_req_bits_in3;
  wire  core_io_fpu_cp_resp_ready;
  wire  core_io_fpu_cp_resp_valid;
  wire [64:0] core_io_fpu_cp_resp_bits_data;
  wire [4:0] core_io_fpu_cp_resp_bits_exc;
  wire  core_io_rocc_cmd_ready;
  wire  core_io_rocc_cmd_valid;
  wire [6:0] core_io_rocc_cmd_bits_inst_funct;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire  core_io_rocc_cmd_bits_inst_xd;
  wire  core_io_rocc_cmd_bits_inst_xs1;
  wire  core_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rd;
  wire [6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire [63:0] core_io_rocc_cmd_bits_rs1;
  wire [63:0] core_io_rocc_cmd_bits_rs2;
  wire  core_io_rocc_resp_ready;
  wire  core_io_rocc_resp_valid;
  wire [4:0] core_io_rocc_resp_bits_rd;
  wire [63:0] core_io_rocc_resp_bits_data;
  wire  core_io_rocc_mem_req_ready;
  wire  core_io_rocc_mem_req_valid;
  wire [39:0] core_io_rocc_mem_req_bits_addr;
  wire [8:0] core_io_rocc_mem_req_bits_tag;
  wire [4:0] core_io_rocc_mem_req_bits_cmd;
  wire [2:0] core_io_rocc_mem_req_bits_typ;
  wire  core_io_rocc_mem_req_bits_phys;
  wire [63:0] core_io_rocc_mem_req_bits_data;
  wire  core_io_rocc_mem_s1_kill;
  wire [63:0] core_io_rocc_mem_s1_data;
  wire  core_io_rocc_mem_s2_nack;
  wire  core_io_rocc_mem_resp_valid;
  wire [39:0] core_io_rocc_mem_resp_bits_addr;
  wire [8:0] core_io_rocc_mem_resp_bits_tag;
  wire [4:0] core_io_rocc_mem_resp_bits_cmd;
  wire [2:0] core_io_rocc_mem_resp_bits_typ;
  wire [63:0] core_io_rocc_mem_resp_bits_data;
  wire  core_io_rocc_mem_resp_bits_replay;
  wire  core_io_rocc_mem_resp_bits_has_data;
  wire [63:0] core_io_rocc_mem_resp_bits_data_word_bypass;
  wire [63:0] core_io_rocc_mem_resp_bits_store_data;
  wire  core_io_rocc_mem_replay_next;
  wire  core_io_rocc_mem_xcpt_ma_ld;
  wire  core_io_rocc_mem_xcpt_ma_st;
  wire  core_io_rocc_mem_xcpt_pf_ld;
  wire  core_io_rocc_mem_xcpt_pf_st;
  wire  core_io_rocc_mem_invalidate_lr;
  wire  core_io_rocc_mem_ordered;
  wire  core_io_rocc_busy;
  wire  core_io_rocc_status_debug;
  wire [1:0] core_io_rocc_status_prv;
  wire  core_io_rocc_status_sd;
  wire [30:0] core_io_rocc_status_zero3;
  wire  core_io_rocc_status_sd_rv32;
  wire [1:0] core_io_rocc_status_zero2;
  wire [4:0] core_io_rocc_status_vm;
  wire [4:0] core_io_rocc_status_zero1;
  wire  core_io_rocc_status_pum;
  wire  core_io_rocc_status_mprv;
  wire [1:0] core_io_rocc_status_xs;
  wire [1:0] core_io_rocc_status_fs;
  wire [1:0] core_io_rocc_status_mpp;
  wire [1:0] core_io_rocc_status_hpp;
  wire  core_io_rocc_status_spp;
  wire  core_io_rocc_status_mpie;
  wire  core_io_rocc_status_hpie;
  wire  core_io_rocc_status_spie;
  wire  core_io_rocc_status_upie;
  wire  core_io_rocc_status_mie;
  wire  core_io_rocc_status_hie;
  wire  core_io_rocc_status_sie;
  wire  core_io_rocc_status_uie;
  wire  core_io_rocc_interrupt;
  wire  core_io_rocc_autl_acquire_ready;
  wire  core_io_rocc_autl_acquire_valid;
  wire [25:0] core_io_rocc_autl_acquire_bits_addr_block;
  wire [1:0] core_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_acquire_bits_addr_beat;
  wire  core_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] core_io_rocc_autl_acquire_bits_a_type;
  wire [11:0] core_io_rocc_autl_acquire_bits_union;
  wire [63:0] core_io_rocc_autl_acquire_bits_data;
  wire  core_io_rocc_autl_grant_ready;
  wire  core_io_rocc_autl_grant_valid;
  wire [2:0] core_io_rocc_autl_grant_bits_addr_beat;
  wire [1:0] core_io_rocc_autl_grant_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_grant_bits_manager_xact_id;
  wire  core_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] core_io_rocc_autl_grant_bits_g_type;
  wire [63:0] core_io_rocc_autl_grant_bits_data;
  wire  core_io_rocc_fpu_req_ready;
  wire  core_io_rocc_fpu_req_valid;
  wire [4:0] core_io_rocc_fpu_req_bits_cmd;
  wire  core_io_rocc_fpu_req_bits_ldst;
  wire  core_io_rocc_fpu_req_bits_wen;
  wire  core_io_rocc_fpu_req_bits_ren1;
  wire  core_io_rocc_fpu_req_bits_ren2;
  wire  core_io_rocc_fpu_req_bits_ren3;
  wire  core_io_rocc_fpu_req_bits_swap12;
  wire  core_io_rocc_fpu_req_bits_swap23;
  wire  core_io_rocc_fpu_req_bits_single;
  wire  core_io_rocc_fpu_req_bits_fromint;
  wire  core_io_rocc_fpu_req_bits_toint;
  wire  core_io_rocc_fpu_req_bits_fastpipe;
  wire  core_io_rocc_fpu_req_bits_fma;
  wire  core_io_rocc_fpu_req_bits_div;
  wire  core_io_rocc_fpu_req_bits_sqrt;
  wire  core_io_rocc_fpu_req_bits_round;
  wire  core_io_rocc_fpu_req_bits_wflags;
  wire [2:0] core_io_rocc_fpu_req_bits_rm;
  wire [1:0] core_io_rocc_fpu_req_bits_typ;
  wire [64:0] core_io_rocc_fpu_req_bits_in1;
  wire [64:0] core_io_rocc_fpu_req_bits_in2;
  wire [64:0] core_io_rocc_fpu_req_bits_in3;
  wire  core_io_rocc_fpu_resp_ready;
  wire  core_io_rocc_fpu_resp_valid;
  wire [64:0] core_io_rocc_fpu_resp_bits_data;
  wire [4:0] core_io_rocc_fpu_resp_bits_exc;
  wire  core_io_rocc_exception;
  wire [11:0] core_io_rocc_csr_waddr;
  wire [63:0] core_io_rocc_csr_wdata;
  wire  core_io_rocc_csr_wen;
  wire  core_io_rocc_host_id;
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_cpu_req_valid;
  wire [39:0] icache_io_cpu_req_bits_pc;
  wire  icache_io_cpu_resp_ready;
  wire  icache_io_cpu_resp_valid;
  wire [39:0] icache_io_cpu_resp_bits_pc;
  wire [31:0] icache_io_cpu_resp_bits_data_0;
  wire  icache_io_cpu_resp_bits_mask;
  wire  icache_io_cpu_resp_bits_xcpt_if;
  wire  icache_io_cpu_btb_resp_valid;
  wire  icache_io_cpu_btb_resp_bits_taken;
  wire  icache_io_cpu_btb_resp_bits_mask;
  wire  icache_io_cpu_btb_resp_bits_bridx;
  wire [38:0] icache_io_cpu_btb_resp_bits_target;
  wire [5:0] icache_io_cpu_btb_resp_bits_entry;
  wire [6:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire  icache_io_cpu_btb_update_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_btb_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_btb_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] icache_io_cpu_btb_update_bits_pc;
  wire [38:0] icache_io_cpu_btb_update_bits_target;
  wire  icache_io_cpu_btb_update_bits_taken;
  wire  icache_io_cpu_btb_update_bits_isJump;
  wire  icache_io_cpu_btb_update_bits_isReturn;
  wire [38:0] icache_io_cpu_btb_update_bits_br_pc;
  wire  icache_io_cpu_bht_update_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_bht_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_bht_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] icache_io_cpu_bht_update_bits_pc;
  wire  icache_io_cpu_bht_update_bits_taken;
  wire  icache_io_cpu_bht_update_bits_mispredict;
  wire  icache_io_cpu_ras_update_valid;
  wire  icache_io_cpu_ras_update_bits_isCall;
  wire  icache_io_cpu_ras_update_bits_isReturn;
  wire [38:0] icache_io_cpu_ras_update_bits_returnAddr;
  wire  icache_io_cpu_ras_update_bits_prediction_valid;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_ras_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_ras_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_value;
  wire  icache_io_cpu_flush_icache;
  wire  icache_io_cpu_flush_tlb;
  wire [39:0] icache_io_cpu_npc;
  wire  icache_io_ptw_req_ready;
  wire  icache_io_ptw_req_valid;
  wire [26:0] icache_io_ptw_req_bits_addr;
  wire [1:0] icache_io_ptw_req_bits_prv;
  wire  icache_io_ptw_req_bits_store;
  wire  icache_io_ptw_req_bits_fetch;
  wire  icache_io_ptw_resp_valid;
  wire [19:0] icache_io_ptw_resp_bits_pte_ppn;
  wire [2:0] icache_io_ptw_resp_bits_pte_reserved_for_software;
  wire  icache_io_ptw_resp_bits_pte_d;
  wire  icache_io_ptw_resp_bits_pte_r;
  wire [3:0] icache_io_ptw_resp_bits_pte_typ;
  wire  icache_io_ptw_resp_bits_pte_v;
  wire [6:0] icache_io_ptw_ptbr_asid;
  wire [37:0] icache_io_ptw_ptbr_ppn;
  wire  icache_io_ptw_invalidate;
  wire  icache_io_ptw_status_debug;
  wire [1:0] icache_io_ptw_status_prv;
  wire  icache_io_ptw_status_sd;
  wire [30:0] icache_io_ptw_status_zero3;
  wire  icache_io_ptw_status_sd_rv32;
  wire [1:0] icache_io_ptw_status_zero2;
  wire [4:0] icache_io_ptw_status_vm;
  wire [4:0] icache_io_ptw_status_zero1;
  wire  icache_io_ptw_status_pum;
  wire  icache_io_ptw_status_mprv;
  wire [1:0] icache_io_ptw_status_xs;
  wire [1:0] icache_io_ptw_status_fs;
  wire [1:0] icache_io_ptw_status_mpp;
  wire [1:0] icache_io_ptw_status_hpp;
  wire  icache_io_ptw_status_spp;
  wire  icache_io_ptw_status_mpie;
  wire  icache_io_ptw_status_hpie;
  wire  icache_io_ptw_status_spie;
  wire  icache_io_ptw_status_upie;
  wire  icache_io_ptw_status_mie;
  wire  icache_io_ptw_status_hie;
  wire  icache_io_ptw_status_sie;
  wire  icache_io_ptw_status_uie;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire [1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [11:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire [1:0] icache_io_mem_grant_bits_client_xact_id;
  wire [2:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  HellaCache_1_clk;
  wire  HellaCache_1_reset;
  wire  HellaCache_1_io_cpu_req_ready;
  wire  HellaCache_1_io_cpu_req_valid;
  wire [39:0] HellaCache_1_io_cpu_req_bits_addr;
  wire [8:0] HellaCache_1_io_cpu_req_bits_tag;
  wire [4:0] HellaCache_1_io_cpu_req_bits_cmd;
  wire [2:0] HellaCache_1_io_cpu_req_bits_typ;
  wire  HellaCache_1_io_cpu_req_bits_phys;
  wire [63:0] HellaCache_1_io_cpu_req_bits_data;
  wire  HellaCache_1_io_cpu_s1_kill;
  wire [63:0] HellaCache_1_io_cpu_s1_data;
  wire  HellaCache_1_io_cpu_s2_nack;
  wire  HellaCache_1_io_cpu_resp_valid;
  wire [39:0] HellaCache_1_io_cpu_resp_bits_addr;
  wire [8:0] HellaCache_1_io_cpu_resp_bits_tag;
  wire [4:0] HellaCache_1_io_cpu_resp_bits_cmd;
  wire [2:0] HellaCache_1_io_cpu_resp_bits_typ;
  wire [63:0] HellaCache_1_io_cpu_resp_bits_data;
  wire  HellaCache_1_io_cpu_resp_bits_replay;
  wire  HellaCache_1_io_cpu_resp_bits_has_data;
  wire [63:0] HellaCache_1_io_cpu_resp_bits_data_word_bypass;
  wire [63:0] HellaCache_1_io_cpu_resp_bits_store_data;
  wire  HellaCache_1_io_cpu_replay_next;
  wire  HellaCache_1_io_cpu_xcpt_ma_ld;
  wire  HellaCache_1_io_cpu_xcpt_ma_st;
  wire  HellaCache_1_io_cpu_xcpt_pf_ld;
  wire  HellaCache_1_io_cpu_xcpt_pf_st;
  wire  HellaCache_1_io_cpu_invalidate_lr;
  wire  HellaCache_1_io_cpu_ordered;
  wire  HellaCache_1_io_ptw_req_ready;
  wire  HellaCache_1_io_ptw_req_valid;
  wire [26:0] HellaCache_1_io_ptw_req_bits_addr;
  wire [1:0] HellaCache_1_io_ptw_req_bits_prv;
  wire  HellaCache_1_io_ptw_req_bits_store;
  wire  HellaCache_1_io_ptw_req_bits_fetch;
  wire  HellaCache_1_io_ptw_resp_valid;
  wire [19:0] HellaCache_1_io_ptw_resp_bits_pte_ppn;
  wire [2:0] HellaCache_1_io_ptw_resp_bits_pte_reserved_for_software;
  wire  HellaCache_1_io_ptw_resp_bits_pte_d;
  wire  HellaCache_1_io_ptw_resp_bits_pte_r;
  wire [3:0] HellaCache_1_io_ptw_resp_bits_pte_typ;
  wire  HellaCache_1_io_ptw_resp_bits_pte_v;
  wire [6:0] HellaCache_1_io_ptw_ptbr_asid;
  wire [37:0] HellaCache_1_io_ptw_ptbr_ppn;
  wire  HellaCache_1_io_ptw_invalidate;
  wire  HellaCache_1_io_ptw_status_debug;
  wire [1:0] HellaCache_1_io_ptw_status_prv;
  wire  HellaCache_1_io_ptw_status_sd;
  wire [30:0] HellaCache_1_io_ptw_status_zero3;
  wire  HellaCache_1_io_ptw_status_sd_rv32;
  wire [1:0] HellaCache_1_io_ptw_status_zero2;
  wire [4:0] HellaCache_1_io_ptw_status_vm;
  wire [4:0] HellaCache_1_io_ptw_status_zero1;
  wire  HellaCache_1_io_ptw_status_pum;
  wire  HellaCache_1_io_ptw_status_mprv;
  wire [1:0] HellaCache_1_io_ptw_status_xs;
  wire [1:0] HellaCache_1_io_ptw_status_fs;
  wire [1:0] HellaCache_1_io_ptw_status_mpp;
  wire [1:0] HellaCache_1_io_ptw_status_hpp;
  wire  HellaCache_1_io_ptw_status_spp;
  wire  HellaCache_1_io_ptw_status_mpie;
  wire  HellaCache_1_io_ptw_status_hpie;
  wire  HellaCache_1_io_ptw_status_spie;
  wire  HellaCache_1_io_ptw_status_upie;
  wire  HellaCache_1_io_ptw_status_mie;
  wire  HellaCache_1_io_ptw_status_hie;
  wire  HellaCache_1_io_ptw_status_sie;
  wire  HellaCache_1_io_ptw_status_uie;
  wire  HellaCache_1_io_mem_acquire_ready;
  wire  HellaCache_1_io_mem_acquire_valid;
  wire [25:0] HellaCache_1_io_mem_acquire_bits_addr_block;
  wire [1:0] HellaCache_1_io_mem_acquire_bits_client_xact_id;
  wire [2:0] HellaCache_1_io_mem_acquire_bits_addr_beat;
  wire  HellaCache_1_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] HellaCache_1_io_mem_acquire_bits_a_type;
  wire [11:0] HellaCache_1_io_mem_acquire_bits_union;
  wire [63:0] HellaCache_1_io_mem_acquire_bits_data;
  wire  HellaCache_1_io_mem_probe_ready;
  wire  HellaCache_1_io_mem_probe_valid;
  wire [25:0] HellaCache_1_io_mem_probe_bits_addr_block;
  wire [1:0] HellaCache_1_io_mem_probe_bits_p_type;
  wire  HellaCache_1_io_mem_release_ready;
  wire  HellaCache_1_io_mem_release_valid;
  wire [2:0] HellaCache_1_io_mem_release_bits_addr_beat;
  wire [25:0] HellaCache_1_io_mem_release_bits_addr_block;
  wire [1:0] HellaCache_1_io_mem_release_bits_client_xact_id;
  wire  HellaCache_1_io_mem_release_bits_voluntary;
  wire [2:0] HellaCache_1_io_mem_release_bits_r_type;
  wire [63:0] HellaCache_1_io_mem_release_bits_data;
  wire  HellaCache_1_io_mem_grant_ready;
  wire  HellaCache_1_io_mem_grant_valid;
  wire [2:0] HellaCache_1_io_mem_grant_bits_addr_beat;
  wire [1:0] HellaCache_1_io_mem_grant_bits_client_xact_id;
  wire [2:0] HellaCache_1_io_mem_grant_bits_manager_xact_id;
  wire  HellaCache_1_io_mem_grant_bits_is_builtin_type;
  wire [3:0] HellaCache_1_io_mem_grant_bits_g_type;
  wire [63:0] HellaCache_1_io_mem_grant_bits_data;
  wire  HellaCache_1_io_mem_grant_bits_manager_id;
  wire  HellaCache_1_io_mem_finish_ready;
  wire  HellaCache_1_io_mem_finish_valid;
  wire [2:0] HellaCache_1_io_mem_finish_bits_manager_xact_id;
  wire  HellaCache_1_io_mem_finish_bits_manager_id;
  wire  uncachedArb_clk;
  wire  uncachedArb_reset;
  wire  uncachedArb_io_in_0_acquire_ready;
  wire  uncachedArb_io_in_0_acquire_valid;
  wire [25:0] uncachedArb_io_in_0_acquire_bits_addr_block;
  wire [1:0] uncachedArb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_addr_beat;
  wire  uncachedArb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_a_type;
  wire [11:0] uncachedArb_io_in_0_acquire_bits_union;
  wire [63:0] uncachedArb_io_in_0_acquire_bits_data;
  wire  uncachedArb_io_in_0_grant_ready;
  wire  uncachedArb_io_in_0_grant_valid;
  wire [2:0] uncachedArb_io_in_0_grant_bits_addr_beat;
  wire [1:0] uncachedArb_io_in_0_grant_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_grant_bits_manager_xact_id;
  wire  uncachedArb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_in_0_grant_bits_g_type;
  wire [63:0] uncachedArb_io_in_0_grant_bits_data;
  wire  uncachedArb_io_out_acquire_ready;
  wire  uncachedArb_io_out_acquire_valid;
  wire [25:0] uncachedArb_io_out_acquire_bits_addr_block;
  wire [1:0] uncachedArb_io_out_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_acquire_bits_addr_beat;
  wire  uncachedArb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_out_acquire_bits_a_type;
  wire [11:0] uncachedArb_io_out_acquire_bits_union;
  wire [63:0] uncachedArb_io_out_acquire_bits_data;
  wire  uncachedArb_io_out_grant_ready;
  wire  uncachedArb_io_out_grant_valid;
  wire [2:0] uncachedArb_io_out_grant_bits_addr_beat;
  wire [1:0] uncachedArb_io_out_grant_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_grant_bits_manager_xact_id;
  wire  uncachedArb_io_out_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_out_grant_bits_g_type;
  wire [63:0] uncachedArb_io_out_grant_bits_data;
  wire  PTW_1_clk;
  wire  PTW_1_reset;
  wire  PTW_1_io_requestor_0_req_ready;
  wire  PTW_1_io_requestor_0_req_valid;
  wire [26:0] PTW_1_io_requestor_0_req_bits_addr;
  wire [1:0] PTW_1_io_requestor_0_req_bits_prv;
  wire  PTW_1_io_requestor_0_req_bits_store;
  wire  PTW_1_io_requestor_0_req_bits_fetch;
  wire  PTW_1_io_requestor_0_resp_valid;
  wire [19:0] PTW_1_io_requestor_0_resp_bits_pte_ppn;
  wire [2:0] PTW_1_io_requestor_0_resp_bits_pte_reserved_for_software;
  wire  PTW_1_io_requestor_0_resp_bits_pte_d;
  wire  PTW_1_io_requestor_0_resp_bits_pte_r;
  wire [3:0] PTW_1_io_requestor_0_resp_bits_pte_typ;
  wire  PTW_1_io_requestor_0_resp_bits_pte_v;
  wire [6:0] PTW_1_io_requestor_0_ptbr_asid;
  wire [37:0] PTW_1_io_requestor_0_ptbr_ppn;
  wire  PTW_1_io_requestor_0_invalidate;
  wire  PTW_1_io_requestor_0_status_debug;
  wire [1:0] PTW_1_io_requestor_0_status_prv;
  wire  PTW_1_io_requestor_0_status_sd;
  wire [30:0] PTW_1_io_requestor_0_status_zero3;
  wire  PTW_1_io_requestor_0_status_sd_rv32;
  wire [1:0] PTW_1_io_requestor_0_status_zero2;
  wire [4:0] PTW_1_io_requestor_0_status_vm;
  wire [4:0] PTW_1_io_requestor_0_status_zero1;
  wire  PTW_1_io_requestor_0_status_pum;
  wire  PTW_1_io_requestor_0_status_mprv;
  wire [1:0] PTW_1_io_requestor_0_status_xs;
  wire [1:0] PTW_1_io_requestor_0_status_fs;
  wire [1:0] PTW_1_io_requestor_0_status_mpp;
  wire [1:0] PTW_1_io_requestor_0_status_hpp;
  wire  PTW_1_io_requestor_0_status_spp;
  wire  PTW_1_io_requestor_0_status_mpie;
  wire  PTW_1_io_requestor_0_status_hpie;
  wire  PTW_1_io_requestor_0_status_spie;
  wire  PTW_1_io_requestor_0_status_upie;
  wire  PTW_1_io_requestor_0_status_mie;
  wire  PTW_1_io_requestor_0_status_hie;
  wire  PTW_1_io_requestor_0_status_sie;
  wire  PTW_1_io_requestor_0_status_uie;
  wire  PTW_1_io_requestor_1_req_ready;
  wire  PTW_1_io_requestor_1_req_valid;
  wire [26:0] PTW_1_io_requestor_1_req_bits_addr;
  wire [1:0] PTW_1_io_requestor_1_req_bits_prv;
  wire  PTW_1_io_requestor_1_req_bits_store;
  wire  PTW_1_io_requestor_1_req_bits_fetch;
  wire  PTW_1_io_requestor_1_resp_valid;
  wire [19:0] PTW_1_io_requestor_1_resp_bits_pte_ppn;
  wire [2:0] PTW_1_io_requestor_1_resp_bits_pte_reserved_for_software;
  wire  PTW_1_io_requestor_1_resp_bits_pte_d;
  wire  PTW_1_io_requestor_1_resp_bits_pte_r;
  wire [3:0] PTW_1_io_requestor_1_resp_bits_pte_typ;
  wire  PTW_1_io_requestor_1_resp_bits_pte_v;
  wire [6:0] PTW_1_io_requestor_1_ptbr_asid;
  wire [37:0] PTW_1_io_requestor_1_ptbr_ppn;
  wire  PTW_1_io_requestor_1_invalidate;
  wire  PTW_1_io_requestor_1_status_debug;
  wire [1:0] PTW_1_io_requestor_1_status_prv;
  wire  PTW_1_io_requestor_1_status_sd;
  wire [30:0] PTW_1_io_requestor_1_status_zero3;
  wire  PTW_1_io_requestor_1_status_sd_rv32;
  wire [1:0] PTW_1_io_requestor_1_status_zero2;
  wire [4:0] PTW_1_io_requestor_1_status_vm;
  wire [4:0] PTW_1_io_requestor_1_status_zero1;
  wire  PTW_1_io_requestor_1_status_pum;
  wire  PTW_1_io_requestor_1_status_mprv;
  wire [1:0] PTW_1_io_requestor_1_status_xs;
  wire [1:0] PTW_1_io_requestor_1_status_fs;
  wire [1:0] PTW_1_io_requestor_1_status_mpp;
  wire [1:0] PTW_1_io_requestor_1_status_hpp;
  wire  PTW_1_io_requestor_1_status_spp;
  wire  PTW_1_io_requestor_1_status_mpie;
  wire  PTW_1_io_requestor_1_status_hpie;
  wire  PTW_1_io_requestor_1_status_spie;
  wire  PTW_1_io_requestor_1_status_upie;
  wire  PTW_1_io_requestor_1_status_mie;
  wire  PTW_1_io_requestor_1_status_hie;
  wire  PTW_1_io_requestor_1_status_sie;
  wire  PTW_1_io_requestor_1_status_uie;
  wire  PTW_1_io_mem_req_ready;
  wire  PTW_1_io_mem_req_valid;
  wire [39:0] PTW_1_io_mem_req_bits_addr;
  wire [8:0] PTW_1_io_mem_req_bits_tag;
  wire [4:0] PTW_1_io_mem_req_bits_cmd;
  wire [2:0] PTW_1_io_mem_req_bits_typ;
  wire  PTW_1_io_mem_req_bits_phys;
  wire [63:0] PTW_1_io_mem_req_bits_data;
  wire  PTW_1_io_mem_s1_kill;
  wire [63:0] PTW_1_io_mem_s1_data;
  wire  PTW_1_io_mem_s2_nack;
  wire  PTW_1_io_mem_resp_valid;
  wire [39:0] PTW_1_io_mem_resp_bits_addr;
  wire [8:0] PTW_1_io_mem_resp_bits_tag;
  wire [4:0] PTW_1_io_mem_resp_bits_cmd;
  wire [2:0] PTW_1_io_mem_resp_bits_typ;
  wire [63:0] PTW_1_io_mem_resp_bits_data;
  wire  PTW_1_io_mem_resp_bits_replay;
  wire  PTW_1_io_mem_resp_bits_has_data;
  wire [63:0] PTW_1_io_mem_resp_bits_data_word_bypass;
  wire [63:0] PTW_1_io_mem_resp_bits_store_data;
  wire  PTW_1_io_mem_replay_next;
  wire  PTW_1_io_mem_xcpt_ma_ld;
  wire  PTW_1_io_mem_xcpt_ma_st;
  wire  PTW_1_io_mem_xcpt_pf_ld;
  wire  PTW_1_io_mem_xcpt_pf_st;
  wire  PTW_1_io_mem_invalidate_lr;
  wire  PTW_1_io_mem_ordered;
  wire [6:0] PTW_1_io_dpath_ptbr_asid;
  wire [37:0] PTW_1_io_dpath_ptbr_ppn;
  wire  PTW_1_io_dpath_invalidate;
  wire  PTW_1_io_dpath_status_debug;
  wire [1:0] PTW_1_io_dpath_status_prv;
  wire  PTW_1_io_dpath_status_sd;
  wire [30:0] PTW_1_io_dpath_status_zero3;
  wire  PTW_1_io_dpath_status_sd_rv32;
  wire [1:0] PTW_1_io_dpath_status_zero2;
  wire [4:0] PTW_1_io_dpath_status_vm;
  wire [4:0] PTW_1_io_dpath_status_zero1;
  wire  PTW_1_io_dpath_status_pum;
  wire  PTW_1_io_dpath_status_mprv;
  wire [1:0] PTW_1_io_dpath_status_xs;
  wire [1:0] PTW_1_io_dpath_status_fs;
  wire [1:0] PTW_1_io_dpath_status_mpp;
  wire [1:0] PTW_1_io_dpath_status_hpp;
  wire  PTW_1_io_dpath_status_spp;
  wire  PTW_1_io_dpath_status_mpie;
  wire  PTW_1_io_dpath_status_hpie;
  wire  PTW_1_io_dpath_status_spie;
  wire  PTW_1_io_dpath_status_upie;
  wire  PTW_1_io_dpath_status_mie;
  wire  PTW_1_io_dpath_status_hie;
  wire  PTW_1_io_dpath_status_sie;
  wire  PTW_1_io_dpath_status_uie;
  wire  dcArb_clk;
  wire  dcArb_reset;
  wire  dcArb_io_requestor_0_req_ready;
  wire  dcArb_io_requestor_0_req_valid;
  wire [39:0] dcArb_io_requestor_0_req_bits_addr;
  wire [8:0] dcArb_io_requestor_0_req_bits_tag;
  wire [4:0] dcArb_io_requestor_0_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_req_bits_typ;
  wire  dcArb_io_requestor_0_req_bits_phys;
  wire [63:0] dcArb_io_requestor_0_req_bits_data;
  wire  dcArb_io_requestor_0_s1_kill;
  wire [63:0] dcArb_io_requestor_0_s1_data;
  wire  dcArb_io_requestor_0_s2_nack;
  wire  dcArb_io_requestor_0_resp_valid;
  wire [39:0] dcArb_io_requestor_0_resp_bits_addr;
  wire [8:0] dcArb_io_requestor_0_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire [63:0] dcArb_io_requestor_0_resp_bits_data;
  wire  dcArb_io_requestor_0_resp_bits_replay;
  wire  dcArb_io_requestor_0_resp_bits_has_data;
  wire [63:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire  dcArb_io_requestor_0_replay_next;
  wire  dcArb_io_requestor_0_xcpt_ma_ld;
  wire  dcArb_io_requestor_0_xcpt_ma_st;
  wire  dcArb_io_requestor_0_xcpt_pf_ld;
  wire  dcArb_io_requestor_0_xcpt_pf_st;
  wire  dcArb_io_requestor_0_invalidate_lr;
  wire  dcArb_io_requestor_0_ordered;
  wire  dcArb_io_requestor_1_req_ready;
  wire  dcArb_io_requestor_1_req_valid;
  wire [39:0] dcArb_io_requestor_1_req_bits_addr;
  wire [8:0] dcArb_io_requestor_1_req_bits_tag;
  wire [4:0] dcArb_io_requestor_1_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_1_req_bits_typ;
  wire  dcArb_io_requestor_1_req_bits_phys;
  wire [63:0] dcArb_io_requestor_1_req_bits_data;
  wire  dcArb_io_requestor_1_s1_kill;
  wire [63:0] dcArb_io_requestor_1_s1_data;
  wire  dcArb_io_requestor_1_s2_nack;
  wire  dcArb_io_requestor_1_resp_valid;
  wire [39:0] dcArb_io_requestor_1_resp_bits_addr;
  wire [8:0] dcArb_io_requestor_1_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire [63:0] dcArb_io_requestor_1_resp_bits_data;
  wire  dcArb_io_requestor_1_resp_bits_replay;
  wire  dcArb_io_requestor_1_resp_bits_has_data;
  wire [63:0] dcArb_io_requestor_1_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire  dcArb_io_requestor_1_replay_next;
  wire  dcArb_io_requestor_1_xcpt_ma_ld;
  wire  dcArb_io_requestor_1_xcpt_ma_st;
  wire  dcArb_io_requestor_1_xcpt_pf_ld;
  wire  dcArb_io_requestor_1_xcpt_pf_st;
  wire  dcArb_io_requestor_1_invalidate_lr;
  wire  dcArb_io_requestor_1_ordered;
  wire  dcArb_io_mem_req_ready;
  wire  dcArb_io_mem_req_valid;
  wire [39:0] dcArb_io_mem_req_bits_addr;
  wire [8:0] dcArb_io_mem_req_bits_tag;
  wire [4:0] dcArb_io_mem_req_bits_cmd;
  wire [2:0] dcArb_io_mem_req_bits_typ;
  wire  dcArb_io_mem_req_bits_phys;
  wire [63:0] dcArb_io_mem_req_bits_data;
  wire  dcArb_io_mem_s1_kill;
  wire [63:0] dcArb_io_mem_s1_data;
  wire  dcArb_io_mem_s2_nack;
  wire  dcArb_io_mem_resp_valid;
  wire [39:0] dcArb_io_mem_resp_bits_addr;
  wire [8:0] dcArb_io_mem_resp_bits_tag;
  wire [4:0] dcArb_io_mem_resp_bits_cmd;
  wire [2:0] dcArb_io_mem_resp_bits_typ;
  wire [63:0] dcArb_io_mem_resp_bits_data;
  wire  dcArb_io_mem_resp_bits_replay;
  wire  dcArb_io_mem_resp_bits_has_data;
  wire [63:0] dcArb_io_mem_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_mem_resp_bits_store_data;
  wire  dcArb_io_mem_replay_next;
  wire  dcArb_io_mem_xcpt_ma_ld;
  wire  dcArb_io_mem_xcpt_ma_st;
  wire  dcArb_io_mem_xcpt_pf_ld;
  wire  dcArb_io_mem_xcpt_pf_st;
  wire  dcArb_io_mem_invalidate_lr;
  wire  dcArb_io_mem_ordered;
  reg  GEN_0;
  reg [31:0] GEN_80;
  reg [4:0] GEN_1;
  reg [31:0] GEN_81;
  reg [63:0] GEN_2;
  reg [63:0] GEN_82;
  reg [63:0] GEN_3;
  reg [63:0] GEN_83;
  reg  GEN_4;
  reg [31:0] GEN_84;
  reg  GEN_5;
  reg [31:0] GEN_85;
  reg  GEN_6;
  reg [31:0] GEN_86;
  reg [4:0] GEN_7;
  reg [31:0] GEN_87;
  reg  GEN_8;
  reg [31:0] GEN_88;
  reg  GEN_9;
  reg [31:0] GEN_89;
  reg  GEN_10;
  reg [31:0] GEN_90;
  reg  GEN_11;
  reg [31:0] GEN_91;
  reg  GEN_12;
  reg [31:0] GEN_92;
  reg  GEN_13;
  reg [31:0] GEN_93;
  reg  GEN_14;
  reg [31:0] GEN_94;
  reg  GEN_15;
  reg [31:0] GEN_95;
  reg  GEN_16;
  reg [31:0] GEN_96;
  reg  GEN_17;
  reg [31:0] GEN_97;
  reg  GEN_18;
  reg [31:0] GEN_98;
  reg  GEN_19;
  reg [31:0] GEN_99;
  reg  GEN_20;
  reg [31:0] GEN_100;
  reg  GEN_21;
  reg [31:0] GEN_101;
  reg  GEN_22;
  reg [31:0] GEN_102;
  reg  GEN_23;
  reg [31:0] GEN_103;
  reg  GEN_24;
  reg [31:0] GEN_104;
  reg  GEN_25;
  reg [31:0] GEN_105;
  reg [4:0] GEN_26;
  reg [31:0] GEN_106;
  reg  GEN_27;
  reg [31:0] GEN_107;
  reg  GEN_28;
  reg [31:0] GEN_108;
  reg [64:0] GEN_29;
  reg [95:0] GEN_109;
  reg [4:0] GEN_30;
  reg [31:0] GEN_110;
  reg  GEN_31;
  reg [31:0] GEN_111;
  reg  GEN_32;
  reg [31:0] GEN_112;
  reg [4:0] GEN_33;
  reg [31:0] GEN_113;
  reg [63:0] GEN_34;
  reg [63:0] GEN_114;
  reg  GEN_35;
  reg [31:0] GEN_115;
  reg [39:0] GEN_36;
  reg [63:0] GEN_116;
  reg [8:0] GEN_37;
  reg [31:0] GEN_117;
  reg [4:0] GEN_38;
  reg [31:0] GEN_118;
  reg [2:0] GEN_39;
  reg [31:0] GEN_119;
  reg  GEN_40;
  reg [31:0] GEN_120;
  reg [63:0] GEN_41;
  reg [63:0] GEN_121;
  reg  GEN_42;
  reg [31:0] GEN_122;
  reg [63:0] GEN_43;
  reg [63:0] GEN_123;
  reg  GEN_44;
  reg [31:0] GEN_124;
  reg  GEN_45;
  reg [31:0] GEN_125;
  reg  GEN_46;
  reg [31:0] GEN_126;
  reg  GEN_47;
  reg [31:0] GEN_127;
  reg [25:0] GEN_48;
  reg [31:0] GEN_128;
  reg [1:0] GEN_49;
  reg [31:0] GEN_129;
  reg [2:0] GEN_50;
  reg [31:0] GEN_130;
  reg  GEN_51;
  reg [31:0] GEN_131;
  reg [2:0] GEN_52;
  reg [31:0] GEN_132;
  reg [11:0] GEN_53;
  reg [31:0] GEN_133;
  reg [63:0] GEN_54;
  reg [63:0] GEN_134;
  reg  GEN_55;
  reg [31:0] GEN_135;
  reg  GEN_56;
  reg [31:0] GEN_136;
  reg [4:0] GEN_57;
  reg [31:0] GEN_137;
  reg  GEN_58;
  reg [31:0] GEN_138;
  reg  GEN_59;
  reg [31:0] GEN_139;
  reg  GEN_60;
  reg [31:0] GEN_140;
  reg  GEN_61;
  reg [31:0] GEN_141;
  reg  GEN_62;
  reg [31:0] GEN_142;
  reg  GEN_63;
  reg [31:0] GEN_143;
  reg  GEN_64;
  reg [31:0] GEN_144;
  reg  GEN_65;
  reg [31:0] GEN_145;
  reg  GEN_66;
  reg [31:0] GEN_146;
  reg  GEN_67;
  reg [31:0] GEN_147;
  reg  GEN_68;
  reg [31:0] GEN_148;
  reg  GEN_69;
  reg [31:0] GEN_149;
  reg  GEN_70;
  reg [31:0] GEN_150;
  reg  GEN_71;
  reg [31:0] GEN_151;
  reg  GEN_72;
  reg [31:0] GEN_152;
  reg  GEN_73;
  reg [31:0] GEN_153;
  reg [2:0] GEN_74;
  reg [31:0] GEN_154;
  reg [1:0] GEN_75;
  reg [31:0] GEN_155;
  reg [64:0] GEN_76;
  reg [95:0] GEN_156;
  reg [64:0] GEN_77;
  reg [95:0] GEN_157;
  reg [64:0] GEN_78;
  reg [95:0] GEN_158;
  reg  GEN_79;
  reg [31:0] GEN_159;
  Rocket core (
    .clk(core_clk),
    .reset(core_reset),
    .io_prci_reset(core_io_prci_reset),
    .io_prci_id(core_io_prci_id),
    .io_prci_interrupts_meip(core_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(core_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(core_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(core_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(core_io_prci_interrupts_msip),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data_0(core_io_imem_resp_bits_data_0),
    .io_imem_resp_bits_mask(core_io_imem_resp_bits_mask),
    .io_imem_resp_bits_xcpt_if(core_io_imem_resp_bits_xcpt_if),
    .io_imem_btb_resp_valid(core_io_imem_btb_resp_valid),
    .io_imem_btb_resp_bits_taken(core_io_imem_btb_resp_bits_taken),
    .io_imem_btb_resp_bits_mask(core_io_imem_btb_resp_bits_mask),
    .io_imem_btb_resp_bits_bridx(core_io_imem_btb_resp_bits_bridx),
    .io_imem_btb_resp_bits_target(core_io_imem_btb_resp_bits_target),
    .io_imem_btb_resp_bits_entry(core_io_imem_btb_resp_bits_entry),
    .io_imem_btb_resp_bits_bht_history(core_io_imem_btb_resp_bits_bht_history),
    .io_imem_btb_resp_bits_bht_value(core_io_imem_btb_resp_bits_bht_value),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_valid(core_io_imem_btb_update_bits_prediction_valid),
    .io_imem_btb_update_bits_prediction_bits_taken(core_io_imem_btb_update_bits_prediction_bits_taken),
    .io_imem_btb_update_bits_prediction_bits_mask(core_io_imem_btb_update_bits_prediction_bits_mask),
    .io_imem_btb_update_bits_prediction_bits_bridx(core_io_imem_btb_update_bits_prediction_bits_bridx),
    .io_imem_btb_update_bits_prediction_bits_target(core_io_imem_btb_update_bits_prediction_bits_target),
    .io_imem_btb_update_bits_prediction_bits_entry(core_io_imem_btb_update_bits_prediction_bits_entry),
    .io_imem_btb_update_bits_prediction_bits_bht_history(core_io_imem_btb_update_bits_prediction_bits_bht_history),
    .io_imem_btb_update_bits_prediction_bits_bht_value(core_io_imem_btb_update_bits_prediction_bits_bht_value),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_target(core_io_imem_btb_update_bits_target),
    .io_imem_btb_update_bits_taken(core_io_imem_btb_update_bits_taken),
    .io_imem_btb_update_bits_isJump(core_io_imem_btb_update_bits_isJump),
    .io_imem_btb_update_bits_isReturn(core_io_imem_btb_update_bits_isReturn),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_valid(core_io_imem_bht_update_bits_prediction_valid),
    .io_imem_bht_update_bits_prediction_bits_taken(core_io_imem_bht_update_bits_prediction_bits_taken),
    .io_imem_bht_update_bits_prediction_bits_mask(core_io_imem_bht_update_bits_prediction_bits_mask),
    .io_imem_bht_update_bits_prediction_bits_bridx(core_io_imem_bht_update_bits_prediction_bits_bridx),
    .io_imem_bht_update_bits_prediction_bits_target(core_io_imem_bht_update_bits_prediction_bits_target),
    .io_imem_bht_update_bits_prediction_bits_entry(core_io_imem_bht_update_bits_prediction_bits_entry),
    .io_imem_bht_update_bits_prediction_bits_bht_history(core_io_imem_bht_update_bits_prediction_bits_bht_history),
    .io_imem_bht_update_bits_prediction_bits_bht_value(core_io_imem_bht_update_bits_prediction_bits_bht_value),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_ras_update_valid(core_io_imem_ras_update_valid),
    .io_imem_ras_update_bits_isCall(core_io_imem_ras_update_bits_isCall),
    .io_imem_ras_update_bits_isReturn(core_io_imem_ras_update_bits_isReturn),
    .io_imem_ras_update_bits_returnAddr(core_io_imem_ras_update_bits_returnAddr),
    .io_imem_ras_update_bits_prediction_valid(core_io_imem_ras_update_bits_prediction_valid),
    .io_imem_ras_update_bits_prediction_bits_taken(core_io_imem_ras_update_bits_prediction_bits_taken),
    .io_imem_ras_update_bits_prediction_bits_mask(core_io_imem_ras_update_bits_prediction_bits_mask),
    .io_imem_ras_update_bits_prediction_bits_bridx(core_io_imem_ras_update_bits_prediction_bits_bridx),
    .io_imem_ras_update_bits_prediction_bits_target(core_io_imem_ras_update_bits_prediction_bits_target),
    .io_imem_ras_update_bits_prediction_bits_entry(core_io_imem_ras_update_bits_prediction_bits_entry),
    .io_imem_ras_update_bits_prediction_bits_bht_history(core_io_imem_ras_update_bits_prediction_bits_bht_history),
    .io_imem_ras_update_bits_prediction_bits_bht_value(core_io_imem_ras_update_bits_prediction_bits_bht_value),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_imem_flush_tlb(core_io_imem_flush_tlb),
    .io_imem_npc(core_io_imem_npc),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_req_bits_phys(core_io_dmem_req_bits_phys),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data(core_io_dmem_s1_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_addr(core_io_dmem_resp_bits_addr),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_cmd(core_io_dmem_resp_bits_cmd),
    .io_dmem_resp_bits_typ(core_io_dmem_resp_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_resp_bits_store_data(core_io_dmem_resp_bits_store_data),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_xcpt_ma_ld(core_io_dmem_xcpt_ma_ld),
    .io_dmem_xcpt_ma_st(core_io_dmem_xcpt_ma_st),
    .io_dmem_xcpt_pf_ld(core_io_dmem_xcpt_pf_ld),
    .io_dmem_xcpt_pf_st(core_io_dmem_xcpt_pf_st),
    .io_dmem_invalidate_lr(core_io_dmem_invalidate_lr),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_ptw_ptbr_asid(core_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(core_io_ptw_invalidate),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_sd(core_io_ptw_status_sd),
    .io_ptw_status_zero3(core_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(core_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(core_io_ptw_status_zero2),
    .io_ptw_status_vm(core_io_ptw_status_vm),
    .io_ptw_status_zero1(core_io_ptw_status_zero1),
    .io_ptw_status_pum(core_io_ptw_status_pum),
    .io_ptw_status_mprv(core_io_ptw_status_mprv),
    .io_ptw_status_xs(core_io_ptw_status_xs),
    .io_ptw_status_fs(core_io_ptw_status_fs),
    .io_ptw_status_mpp(core_io_ptw_status_mpp),
    .io_ptw_status_hpp(core_io_ptw_status_hpp),
    .io_ptw_status_spp(core_io_ptw_status_spp),
    .io_ptw_status_mpie(core_io_ptw_status_mpie),
    .io_ptw_status_hpie(core_io_ptw_status_hpie),
    .io_ptw_status_spie(core_io_ptw_status_spie),
    .io_ptw_status_upie(core_io_ptw_status_upie),
    .io_ptw_status_mie(core_io_ptw_status_mie),
    .io_ptw_status_hie(core_io_ptw_status_hie),
    .io_ptw_status_sie(core_io_ptw_status_sie),
    .io_ptw_status_uie(core_io_ptw_status_uie),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_cmd(core_io_fpu_dec_cmd),
    .io_fpu_dec_ldst(core_io_fpu_dec_ldst),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_dec_swap12(core_io_fpu_dec_swap12),
    .io_fpu_dec_swap23(core_io_fpu_dec_swap23),
    .io_fpu_dec_single(core_io_fpu_dec_single),
    .io_fpu_dec_fromint(core_io_fpu_dec_fromint),
    .io_fpu_dec_toint(core_io_fpu_dec_toint),
    .io_fpu_dec_fastpipe(core_io_fpu_dec_fastpipe),
    .io_fpu_dec_fma(core_io_fpu_dec_fma),
    .io_fpu_dec_div(core_io_fpu_dec_div),
    .io_fpu_dec_sqrt(core_io_fpu_dec_sqrt),
    .io_fpu_dec_round(core_io_fpu_dec_round),
    .io_fpu_dec_wflags(core_io_fpu_dec_wflags),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_fpu_cp_req_ready(core_io_fpu_cp_req_ready),
    .io_fpu_cp_req_valid(core_io_fpu_cp_req_valid),
    .io_fpu_cp_req_bits_cmd(core_io_fpu_cp_req_bits_cmd),
    .io_fpu_cp_req_bits_ldst(core_io_fpu_cp_req_bits_ldst),
    .io_fpu_cp_req_bits_wen(core_io_fpu_cp_req_bits_wen),
    .io_fpu_cp_req_bits_ren1(core_io_fpu_cp_req_bits_ren1),
    .io_fpu_cp_req_bits_ren2(core_io_fpu_cp_req_bits_ren2),
    .io_fpu_cp_req_bits_ren3(core_io_fpu_cp_req_bits_ren3),
    .io_fpu_cp_req_bits_swap12(core_io_fpu_cp_req_bits_swap12),
    .io_fpu_cp_req_bits_swap23(core_io_fpu_cp_req_bits_swap23),
    .io_fpu_cp_req_bits_single(core_io_fpu_cp_req_bits_single),
    .io_fpu_cp_req_bits_fromint(core_io_fpu_cp_req_bits_fromint),
    .io_fpu_cp_req_bits_toint(core_io_fpu_cp_req_bits_toint),
    .io_fpu_cp_req_bits_fastpipe(core_io_fpu_cp_req_bits_fastpipe),
    .io_fpu_cp_req_bits_fma(core_io_fpu_cp_req_bits_fma),
    .io_fpu_cp_req_bits_div(core_io_fpu_cp_req_bits_div),
    .io_fpu_cp_req_bits_sqrt(core_io_fpu_cp_req_bits_sqrt),
    .io_fpu_cp_req_bits_round(core_io_fpu_cp_req_bits_round),
    .io_fpu_cp_req_bits_wflags(core_io_fpu_cp_req_bits_wflags),
    .io_fpu_cp_req_bits_rm(core_io_fpu_cp_req_bits_rm),
    .io_fpu_cp_req_bits_typ(core_io_fpu_cp_req_bits_typ),
    .io_fpu_cp_req_bits_in1(core_io_fpu_cp_req_bits_in1),
    .io_fpu_cp_req_bits_in2(core_io_fpu_cp_req_bits_in2),
    .io_fpu_cp_req_bits_in3(core_io_fpu_cp_req_bits_in3),
    .io_fpu_cp_resp_ready(core_io_fpu_cp_resp_ready),
    .io_fpu_cp_resp_valid(core_io_fpu_cp_resp_valid),
    .io_fpu_cp_resp_bits_data(core_io_fpu_cp_resp_bits_data),
    .io_fpu_cp_resp_bits_exc(core_io_fpu_cp_resp_bits_exc),
    .io_rocc_cmd_ready(core_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(core_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(core_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(core_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(core_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(core_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(core_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(core_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(core_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(core_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(core_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(core_io_rocc_cmd_bits_rs2),
    .io_rocc_resp_ready(core_io_rocc_resp_ready),
    .io_rocc_resp_valid(core_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(core_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(core_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(core_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(core_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(core_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(core_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(core_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(core_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(core_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(core_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(core_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(core_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(core_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(core_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(core_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(core_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(core_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(core_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(core_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(core_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(core_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(core_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(core_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(core_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(core_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(core_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(core_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(core_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(core_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(core_io_rocc_mem_ordered),
    .io_rocc_busy(core_io_rocc_busy),
    .io_rocc_status_debug(core_io_rocc_status_debug),
    .io_rocc_status_prv(core_io_rocc_status_prv),
    .io_rocc_status_sd(core_io_rocc_status_sd),
    .io_rocc_status_zero3(core_io_rocc_status_zero3),
    .io_rocc_status_sd_rv32(core_io_rocc_status_sd_rv32),
    .io_rocc_status_zero2(core_io_rocc_status_zero2),
    .io_rocc_status_vm(core_io_rocc_status_vm),
    .io_rocc_status_zero1(core_io_rocc_status_zero1),
    .io_rocc_status_pum(core_io_rocc_status_pum),
    .io_rocc_status_mprv(core_io_rocc_status_mprv),
    .io_rocc_status_xs(core_io_rocc_status_xs),
    .io_rocc_status_fs(core_io_rocc_status_fs),
    .io_rocc_status_mpp(core_io_rocc_status_mpp),
    .io_rocc_status_hpp(core_io_rocc_status_hpp),
    .io_rocc_status_spp(core_io_rocc_status_spp),
    .io_rocc_status_mpie(core_io_rocc_status_mpie),
    .io_rocc_status_hpie(core_io_rocc_status_hpie),
    .io_rocc_status_spie(core_io_rocc_status_spie),
    .io_rocc_status_upie(core_io_rocc_status_upie),
    .io_rocc_status_mie(core_io_rocc_status_mie),
    .io_rocc_status_hie(core_io_rocc_status_hie),
    .io_rocc_status_sie(core_io_rocc_status_sie),
    .io_rocc_status_uie(core_io_rocc_status_uie),
    .io_rocc_interrupt(core_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(core_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(core_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(core_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(core_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(core_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(core_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(core_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(core_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(core_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(core_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(core_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(core_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(core_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(core_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(core_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(core_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(core_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(core_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(core_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(core_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(core_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(core_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(core_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(core_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(core_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(core_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(core_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(core_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(core_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(core_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(core_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(core_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(core_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(core_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(core_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(core_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(core_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(core_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(core_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(core_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(core_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(core_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(core_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(core_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(core_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(core_io_rocc_exception),
    .io_rocc_csr_waddr(core_io_rocc_csr_waddr),
    .io_rocc_csr_wdata(core_io_rocc_csr_wdata),
    .io_rocc_csr_wen(core_io_rocc_csr_wen),
    .io_rocc_host_id(core_io_rocc_host_id)
  );
  Frontend icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_cpu_req_valid(icache_io_cpu_req_valid),
    .io_cpu_req_bits_pc(icache_io_cpu_req_bits_pc),
    .io_cpu_resp_ready(icache_io_cpu_resp_ready),
    .io_cpu_resp_valid(icache_io_cpu_resp_valid),
    .io_cpu_resp_bits_pc(icache_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data_0(icache_io_cpu_resp_bits_data_0),
    .io_cpu_resp_bits_mask(icache_io_cpu_resp_bits_mask),
    .io_cpu_resp_bits_xcpt_if(icache_io_cpu_resp_bits_xcpt_if),
    .io_cpu_btb_resp_valid(icache_io_cpu_btb_resp_valid),
    .io_cpu_btb_resp_bits_taken(icache_io_cpu_btb_resp_bits_taken),
    .io_cpu_btb_resp_bits_mask(icache_io_cpu_btb_resp_bits_mask),
    .io_cpu_btb_resp_bits_bridx(icache_io_cpu_btb_resp_bits_bridx),
    .io_cpu_btb_resp_bits_target(icache_io_cpu_btb_resp_bits_target),
    .io_cpu_btb_resp_bits_entry(icache_io_cpu_btb_resp_bits_entry),
    .io_cpu_btb_resp_bits_bht_history(icache_io_cpu_btb_resp_bits_bht_history),
    .io_cpu_btb_resp_bits_bht_value(icache_io_cpu_btb_resp_bits_bht_value),
    .io_cpu_btb_update_valid(icache_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_valid(icache_io_cpu_btb_update_bits_prediction_valid),
    .io_cpu_btb_update_bits_prediction_bits_taken(icache_io_cpu_btb_update_bits_prediction_bits_taken),
    .io_cpu_btb_update_bits_prediction_bits_mask(icache_io_cpu_btb_update_bits_prediction_bits_mask),
    .io_cpu_btb_update_bits_prediction_bits_bridx(icache_io_cpu_btb_update_bits_prediction_bits_bridx),
    .io_cpu_btb_update_bits_prediction_bits_target(icache_io_cpu_btb_update_bits_prediction_bits_target),
    .io_cpu_btb_update_bits_prediction_bits_entry(icache_io_cpu_btb_update_bits_prediction_bits_entry),
    .io_cpu_btb_update_bits_prediction_bits_bht_history(icache_io_cpu_btb_update_bits_prediction_bits_bht_history),
    .io_cpu_btb_update_bits_prediction_bits_bht_value(icache_io_cpu_btb_update_bits_prediction_bits_bht_value),
    .io_cpu_btb_update_bits_pc(icache_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_target(icache_io_cpu_btb_update_bits_target),
    .io_cpu_btb_update_bits_taken(icache_io_cpu_btb_update_bits_taken),
    .io_cpu_btb_update_bits_isJump(icache_io_cpu_btb_update_bits_isJump),
    .io_cpu_btb_update_bits_isReturn(icache_io_cpu_btb_update_bits_isReturn),
    .io_cpu_btb_update_bits_br_pc(icache_io_cpu_btb_update_bits_br_pc),
    .io_cpu_bht_update_valid(icache_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_valid(icache_io_cpu_bht_update_bits_prediction_valid),
    .io_cpu_bht_update_bits_prediction_bits_taken(icache_io_cpu_bht_update_bits_prediction_bits_taken),
    .io_cpu_bht_update_bits_prediction_bits_mask(icache_io_cpu_bht_update_bits_prediction_bits_mask),
    .io_cpu_bht_update_bits_prediction_bits_bridx(icache_io_cpu_bht_update_bits_prediction_bits_bridx),
    .io_cpu_bht_update_bits_prediction_bits_target(icache_io_cpu_bht_update_bits_prediction_bits_target),
    .io_cpu_bht_update_bits_prediction_bits_entry(icache_io_cpu_bht_update_bits_prediction_bits_entry),
    .io_cpu_bht_update_bits_prediction_bits_bht_history(icache_io_cpu_bht_update_bits_prediction_bits_bht_history),
    .io_cpu_bht_update_bits_prediction_bits_bht_value(icache_io_cpu_bht_update_bits_prediction_bits_bht_value),
    .io_cpu_bht_update_bits_pc(icache_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_taken(icache_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(icache_io_cpu_bht_update_bits_mispredict),
    .io_cpu_ras_update_valid(icache_io_cpu_ras_update_valid),
    .io_cpu_ras_update_bits_isCall(icache_io_cpu_ras_update_bits_isCall),
    .io_cpu_ras_update_bits_isReturn(icache_io_cpu_ras_update_bits_isReturn),
    .io_cpu_ras_update_bits_returnAddr(icache_io_cpu_ras_update_bits_returnAddr),
    .io_cpu_ras_update_bits_prediction_valid(icache_io_cpu_ras_update_bits_prediction_valid),
    .io_cpu_ras_update_bits_prediction_bits_taken(icache_io_cpu_ras_update_bits_prediction_bits_taken),
    .io_cpu_ras_update_bits_prediction_bits_mask(icache_io_cpu_ras_update_bits_prediction_bits_mask),
    .io_cpu_ras_update_bits_prediction_bits_bridx(icache_io_cpu_ras_update_bits_prediction_bits_bridx),
    .io_cpu_ras_update_bits_prediction_bits_target(icache_io_cpu_ras_update_bits_prediction_bits_target),
    .io_cpu_ras_update_bits_prediction_bits_entry(icache_io_cpu_ras_update_bits_prediction_bits_entry),
    .io_cpu_ras_update_bits_prediction_bits_bht_history(icache_io_cpu_ras_update_bits_prediction_bits_bht_history),
    .io_cpu_ras_update_bits_prediction_bits_bht_value(icache_io_cpu_ras_update_bits_prediction_bits_bht_value),
    .io_cpu_flush_icache(icache_io_cpu_flush_icache),
    .io_cpu_flush_tlb(icache_io_cpu_flush_tlb),
    .io_cpu_npc(icache_io_cpu_npc),
    .io_ptw_req_ready(icache_io_ptw_req_ready),
    .io_ptw_req_valid(icache_io_ptw_req_valid),
    .io_ptw_req_bits_addr(icache_io_ptw_req_bits_addr),
    .io_ptw_req_bits_prv(icache_io_ptw_req_bits_prv),
    .io_ptw_req_bits_store(icache_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(icache_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(icache_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_ppn(icache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(icache_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(icache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_r(icache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_typ(icache_io_ptw_resp_bits_pte_typ),
    .io_ptw_resp_bits_pte_v(icache_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(icache_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(icache_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(icache_io_ptw_invalidate),
    .io_ptw_status_debug(icache_io_ptw_status_debug),
    .io_ptw_status_prv(icache_io_ptw_status_prv),
    .io_ptw_status_sd(icache_io_ptw_status_sd),
    .io_ptw_status_zero3(icache_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(icache_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(icache_io_ptw_status_zero2),
    .io_ptw_status_vm(icache_io_ptw_status_vm),
    .io_ptw_status_zero1(icache_io_ptw_status_zero1),
    .io_ptw_status_pum(icache_io_ptw_status_pum),
    .io_ptw_status_mprv(icache_io_ptw_status_mprv),
    .io_ptw_status_xs(icache_io_ptw_status_xs),
    .io_ptw_status_fs(icache_io_ptw_status_fs),
    .io_ptw_status_mpp(icache_io_ptw_status_mpp),
    .io_ptw_status_hpp(icache_io_ptw_status_hpp),
    .io_ptw_status_spp(icache_io_ptw_status_spp),
    .io_ptw_status_mpie(icache_io_ptw_status_mpie),
    .io_ptw_status_hpie(icache_io_ptw_status_hpie),
    .io_ptw_status_spie(icache_io_ptw_status_spie),
    .io_ptw_status_upie(icache_io_ptw_status_upie),
    .io_ptw_status_mie(icache_io_ptw_status_mie),
    .io_ptw_status_hie(icache_io_ptw_status_hie),
    .io_ptw_status_sie(icache_io_ptw_status_sie),
    .io_ptw_status_uie(icache_io_ptw_status_uie),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  HellaCache HellaCache_1 (
    .clk(HellaCache_1_clk),
    .reset(HellaCache_1_reset),
    .io_cpu_req_ready(HellaCache_1_io_cpu_req_ready),
    .io_cpu_req_valid(HellaCache_1_io_cpu_req_valid),
    .io_cpu_req_bits_addr(HellaCache_1_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(HellaCache_1_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(HellaCache_1_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(HellaCache_1_io_cpu_req_bits_typ),
    .io_cpu_req_bits_phys(HellaCache_1_io_cpu_req_bits_phys),
    .io_cpu_req_bits_data(HellaCache_1_io_cpu_req_bits_data),
    .io_cpu_s1_kill(HellaCache_1_io_cpu_s1_kill),
    .io_cpu_s1_data(HellaCache_1_io_cpu_s1_data),
    .io_cpu_s2_nack(HellaCache_1_io_cpu_s2_nack),
    .io_cpu_resp_valid(HellaCache_1_io_cpu_resp_valid),
    .io_cpu_resp_bits_addr(HellaCache_1_io_cpu_resp_bits_addr),
    .io_cpu_resp_bits_tag(HellaCache_1_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_cmd(HellaCache_1_io_cpu_resp_bits_cmd),
    .io_cpu_resp_bits_typ(HellaCache_1_io_cpu_resp_bits_typ),
    .io_cpu_resp_bits_data(HellaCache_1_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(HellaCache_1_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(HellaCache_1_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(HellaCache_1_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_resp_bits_store_data(HellaCache_1_io_cpu_resp_bits_store_data),
    .io_cpu_replay_next(HellaCache_1_io_cpu_replay_next),
    .io_cpu_xcpt_ma_ld(HellaCache_1_io_cpu_xcpt_ma_ld),
    .io_cpu_xcpt_ma_st(HellaCache_1_io_cpu_xcpt_ma_st),
    .io_cpu_xcpt_pf_ld(HellaCache_1_io_cpu_xcpt_pf_ld),
    .io_cpu_xcpt_pf_st(HellaCache_1_io_cpu_xcpt_pf_st),
    .io_cpu_invalidate_lr(HellaCache_1_io_cpu_invalidate_lr),
    .io_cpu_ordered(HellaCache_1_io_cpu_ordered),
    .io_ptw_req_ready(HellaCache_1_io_ptw_req_ready),
    .io_ptw_req_valid(HellaCache_1_io_ptw_req_valid),
    .io_ptw_req_bits_addr(HellaCache_1_io_ptw_req_bits_addr),
    .io_ptw_req_bits_prv(HellaCache_1_io_ptw_req_bits_prv),
    .io_ptw_req_bits_store(HellaCache_1_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(HellaCache_1_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(HellaCache_1_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_ppn(HellaCache_1_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(HellaCache_1_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(HellaCache_1_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_r(HellaCache_1_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_typ(HellaCache_1_io_ptw_resp_bits_pte_typ),
    .io_ptw_resp_bits_pte_v(HellaCache_1_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(HellaCache_1_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(HellaCache_1_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(HellaCache_1_io_ptw_invalidate),
    .io_ptw_status_debug(HellaCache_1_io_ptw_status_debug),
    .io_ptw_status_prv(HellaCache_1_io_ptw_status_prv),
    .io_ptw_status_sd(HellaCache_1_io_ptw_status_sd),
    .io_ptw_status_zero3(HellaCache_1_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(HellaCache_1_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(HellaCache_1_io_ptw_status_zero2),
    .io_ptw_status_vm(HellaCache_1_io_ptw_status_vm),
    .io_ptw_status_zero1(HellaCache_1_io_ptw_status_zero1),
    .io_ptw_status_pum(HellaCache_1_io_ptw_status_pum),
    .io_ptw_status_mprv(HellaCache_1_io_ptw_status_mprv),
    .io_ptw_status_xs(HellaCache_1_io_ptw_status_xs),
    .io_ptw_status_fs(HellaCache_1_io_ptw_status_fs),
    .io_ptw_status_mpp(HellaCache_1_io_ptw_status_mpp),
    .io_ptw_status_hpp(HellaCache_1_io_ptw_status_hpp),
    .io_ptw_status_spp(HellaCache_1_io_ptw_status_spp),
    .io_ptw_status_mpie(HellaCache_1_io_ptw_status_mpie),
    .io_ptw_status_hpie(HellaCache_1_io_ptw_status_hpie),
    .io_ptw_status_spie(HellaCache_1_io_ptw_status_spie),
    .io_ptw_status_upie(HellaCache_1_io_ptw_status_upie),
    .io_ptw_status_mie(HellaCache_1_io_ptw_status_mie),
    .io_ptw_status_hie(HellaCache_1_io_ptw_status_hie),
    .io_ptw_status_sie(HellaCache_1_io_ptw_status_sie),
    .io_ptw_status_uie(HellaCache_1_io_ptw_status_uie),
    .io_mem_acquire_ready(HellaCache_1_io_mem_acquire_ready),
    .io_mem_acquire_valid(HellaCache_1_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(HellaCache_1_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(HellaCache_1_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(HellaCache_1_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(HellaCache_1_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(HellaCache_1_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(HellaCache_1_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(HellaCache_1_io_mem_acquire_bits_data),
    .io_mem_probe_ready(HellaCache_1_io_mem_probe_ready),
    .io_mem_probe_valid(HellaCache_1_io_mem_probe_valid),
    .io_mem_probe_bits_addr_block(HellaCache_1_io_mem_probe_bits_addr_block),
    .io_mem_probe_bits_p_type(HellaCache_1_io_mem_probe_bits_p_type),
    .io_mem_release_ready(HellaCache_1_io_mem_release_ready),
    .io_mem_release_valid(HellaCache_1_io_mem_release_valid),
    .io_mem_release_bits_addr_beat(HellaCache_1_io_mem_release_bits_addr_beat),
    .io_mem_release_bits_addr_block(HellaCache_1_io_mem_release_bits_addr_block),
    .io_mem_release_bits_client_xact_id(HellaCache_1_io_mem_release_bits_client_xact_id),
    .io_mem_release_bits_voluntary(HellaCache_1_io_mem_release_bits_voluntary),
    .io_mem_release_bits_r_type(HellaCache_1_io_mem_release_bits_r_type),
    .io_mem_release_bits_data(HellaCache_1_io_mem_release_bits_data),
    .io_mem_grant_ready(HellaCache_1_io_mem_grant_ready),
    .io_mem_grant_valid(HellaCache_1_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(HellaCache_1_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(HellaCache_1_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(HellaCache_1_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(HellaCache_1_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(HellaCache_1_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(HellaCache_1_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(HellaCache_1_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(HellaCache_1_io_mem_finish_ready),
    .io_mem_finish_valid(HellaCache_1_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(HellaCache_1_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(HellaCache_1_io_mem_finish_bits_manager_id)
  );
  ClientUncachedTileLinkIOArbiter uncachedArb (
    .clk(uncachedArb_clk),
    .reset(uncachedArb_reset),
    .io_in_0_acquire_ready(uncachedArb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(uncachedArb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(uncachedArb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(uncachedArb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(uncachedArb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(uncachedArb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(uncachedArb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(uncachedArb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(uncachedArb_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(uncachedArb_io_in_0_grant_ready),
    .io_in_0_grant_valid(uncachedArb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(uncachedArb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(uncachedArb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(uncachedArb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(uncachedArb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(uncachedArb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(uncachedArb_io_in_0_grant_bits_data),
    .io_out_acquire_ready(uncachedArb_io_out_acquire_ready),
    .io_out_acquire_valid(uncachedArb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(uncachedArb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(uncachedArb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(uncachedArb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(uncachedArb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(uncachedArb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(uncachedArb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(uncachedArb_io_out_acquire_bits_data),
    .io_out_grant_ready(uncachedArb_io_out_grant_ready),
    .io_out_grant_valid(uncachedArb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(uncachedArb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(uncachedArb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(uncachedArb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(uncachedArb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(uncachedArb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(uncachedArb_io_out_grant_bits_data)
  );
  PTW PTW_1 (
    .clk(PTW_1_clk),
    .reset(PTW_1_reset),
    .io_requestor_0_req_ready(PTW_1_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(PTW_1_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(PTW_1_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_prv(PTW_1_io_requestor_0_req_bits_prv),
    .io_requestor_0_req_bits_store(PTW_1_io_requestor_0_req_bits_store),
    .io_requestor_0_req_bits_fetch(PTW_1_io_requestor_0_req_bits_fetch),
    .io_requestor_0_resp_valid(PTW_1_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_pte_ppn(PTW_1_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_reserved_for_software(PTW_1_io_requestor_0_resp_bits_pte_reserved_for_software),
    .io_requestor_0_resp_bits_pte_d(PTW_1_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_r(PTW_1_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_typ(PTW_1_io_requestor_0_resp_bits_pte_typ),
    .io_requestor_0_resp_bits_pte_v(PTW_1_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_ptbr_asid(PTW_1_io_requestor_0_ptbr_asid),
    .io_requestor_0_ptbr_ppn(PTW_1_io_requestor_0_ptbr_ppn),
    .io_requestor_0_invalidate(PTW_1_io_requestor_0_invalidate),
    .io_requestor_0_status_debug(PTW_1_io_requestor_0_status_debug),
    .io_requestor_0_status_prv(PTW_1_io_requestor_0_status_prv),
    .io_requestor_0_status_sd(PTW_1_io_requestor_0_status_sd),
    .io_requestor_0_status_zero3(PTW_1_io_requestor_0_status_zero3),
    .io_requestor_0_status_sd_rv32(PTW_1_io_requestor_0_status_sd_rv32),
    .io_requestor_0_status_zero2(PTW_1_io_requestor_0_status_zero2),
    .io_requestor_0_status_vm(PTW_1_io_requestor_0_status_vm),
    .io_requestor_0_status_zero1(PTW_1_io_requestor_0_status_zero1),
    .io_requestor_0_status_pum(PTW_1_io_requestor_0_status_pum),
    .io_requestor_0_status_mprv(PTW_1_io_requestor_0_status_mprv),
    .io_requestor_0_status_xs(PTW_1_io_requestor_0_status_xs),
    .io_requestor_0_status_fs(PTW_1_io_requestor_0_status_fs),
    .io_requestor_0_status_mpp(PTW_1_io_requestor_0_status_mpp),
    .io_requestor_0_status_hpp(PTW_1_io_requestor_0_status_hpp),
    .io_requestor_0_status_spp(PTW_1_io_requestor_0_status_spp),
    .io_requestor_0_status_mpie(PTW_1_io_requestor_0_status_mpie),
    .io_requestor_0_status_hpie(PTW_1_io_requestor_0_status_hpie),
    .io_requestor_0_status_spie(PTW_1_io_requestor_0_status_spie),
    .io_requestor_0_status_upie(PTW_1_io_requestor_0_status_upie),
    .io_requestor_0_status_mie(PTW_1_io_requestor_0_status_mie),
    .io_requestor_0_status_hie(PTW_1_io_requestor_0_status_hie),
    .io_requestor_0_status_sie(PTW_1_io_requestor_0_status_sie),
    .io_requestor_0_status_uie(PTW_1_io_requestor_0_status_uie),
    .io_requestor_1_req_ready(PTW_1_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(PTW_1_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(PTW_1_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_prv(PTW_1_io_requestor_1_req_bits_prv),
    .io_requestor_1_req_bits_store(PTW_1_io_requestor_1_req_bits_store),
    .io_requestor_1_req_bits_fetch(PTW_1_io_requestor_1_req_bits_fetch),
    .io_requestor_1_resp_valid(PTW_1_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_pte_ppn(PTW_1_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_reserved_for_software(PTW_1_io_requestor_1_resp_bits_pte_reserved_for_software),
    .io_requestor_1_resp_bits_pte_d(PTW_1_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_r(PTW_1_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_typ(PTW_1_io_requestor_1_resp_bits_pte_typ),
    .io_requestor_1_resp_bits_pte_v(PTW_1_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_ptbr_asid(PTW_1_io_requestor_1_ptbr_asid),
    .io_requestor_1_ptbr_ppn(PTW_1_io_requestor_1_ptbr_ppn),
    .io_requestor_1_invalidate(PTW_1_io_requestor_1_invalidate),
    .io_requestor_1_status_debug(PTW_1_io_requestor_1_status_debug),
    .io_requestor_1_status_prv(PTW_1_io_requestor_1_status_prv),
    .io_requestor_1_status_sd(PTW_1_io_requestor_1_status_sd),
    .io_requestor_1_status_zero3(PTW_1_io_requestor_1_status_zero3),
    .io_requestor_1_status_sd_rv32(PTW_1_io_requestor_1_status_sd_rv32),
    .io_requestor_1_status_zero2(PTW_1_io_requestor_1_status_zero2),
    .io_requestor_1_status_vm(PTW_1_io_requestor_1_status_vm),
    .io_requestor_1_status_zero1(PTW_1_io_requestor_1_status_zero1),
    .io_requestor_1_status_pum(PTW_1_io_requestor_1_status_pum),
    .io_requestor_1_status_mprv(PTW_1_io_requestor_1_status_mprv),
    .io_requestor_1_status_xs(PTW_1_io_requestor_1_status_xs),
    .io_requestor_1_status_fs(PTW_1_io_requestor_1_status_fs),
    .io_requestor_1_status_mpp(PTW_1_io_requestor_1_status_mpp),
    .io_requestor_1_status_hpp(PTW_1_io_requestor_1_status_hpp),
    .io_requestor_1_status_spp(PTW_1_io_requestor_1_status_spp),
    .io_requestor_1_status_mpie(PTW_1_io_requestor_1_status_mpie),
    .io_requestor_1_status_hpie(PTW_1_io_requestor_1_status_hpie),
    .io_requestor_1_status_spie(PTW_1_io_requestor_1_status_spie),
    .io_requestor_1_status_upie(PTW_1_io_requestor_1_status_upie),
    .io_requestor_1_status_mie(PTW_1_io_requestor_1_status_mie),
    .io_requestor_1_status_hie(PTW_1_io_requestor_1_status_hie),
    .io_requestor_1_status_sie(PTW_1_io_requestor_1_status_sie),
    .io_requestor_1_status_uie(PTW_1_io_requestor_1_status_uie),
    .io_mem_req_ready(PTW_1_io_mem_req_ready),
    .io_mem_req_valid(PTW_1_io_mem_req_valid),
    .io_mem_req_bits_addr(PTW_1_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(PTW_1_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(PTW_1_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(PTW_1_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(PTW_1_io_mem_req_bits_phys),
    .io_mem_req_bits_data(PTW_1_io_mem_req_bits_data),
    .io_mem_s1_kill(PTW_1_io_mem_s1_kill),
    .io_mem_s1_data(PTW_1_io_mem_s1_data),
    .io_mem_s2_nack(PTW_1_io_mem_s2_nack),
    .io_mem_resp_valid(PTW_1_io_mem_resp_valid),
    .io_mem_resp_bits_addr(PTW_1_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(PTW_1_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(PTW_1_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(PTW_1_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(PTW_1_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(PTW_1_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(PTW_1_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(PTW_1_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(PTW_1_io_mem_resp_bits_store_data),
    .io_mem_replay_next(PTW_1_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(PTW_1_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(PTW_1_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(PTW_1_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(PTW_1_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(PTW_1_io_mem_invalidate_lr),
    .io_mem_ordered(PTW_1_io_mem_ordered),
    .io_dpath_ptbr_asid(PTW_1_io_dpath_ptbr_asid),
    .io_dpath_ptbr_ppn(PTW_1_io_dpath_ptbr_ppn),
    .io_dpath_invalidate(PTW_1_io_dpath_invalidate),
    .io_dpath_status_debug(PTW_1_io_dpath_status_debug),
    .io_dpath_status_prv(PTW_1_io_dpath_status_prv),
    .io_dpath_status_sd(PTW_1_io_dpath_status_sd),
    .io_dpath_status_zero3(PTW_1_io_dpath_status_zero3),
    .io_dpath_status_sd_rv32(PTW_1_io_dpath_status_sd_rv32),
    .io_dpath_status_zero2(PTW_1_io_dpath_status_zero2),
    .io_dpath_status_vm(PTW_1_io_dpath_status_vm),
    .io_dpath_status_zero1(PTW_1_io_dpath_status_zero1),
    .io_dpath_status_pum(PTW_1_io_dpath_status_pum),
    .io_dpath_status_mprv(PTW_1_io_dpath_status_mprv),
    .io_dpath_status_xs(PTW_1_io_dpath_status_xs),
    .io_dpath_status_fs(PTW_1_io_dpath_status_fs),
    .io_dpath_status_mpp(PTW_1_io_dpath_status_mpp),
    .io_dpath_status_hpp(PTW_1_io_dpath_status_hpp),
    .io_dpath_status_spp(PTW_1_io_dpath_status_spp),
    .io_dpath_status_mpie(PTW_1_io_dpath_status_mpie),
    .io_dpath_status_hpie(PTW_1_io_dpath_status_hpie),
    .io_dpath_status_spie(PTW_1_io_dpath_status_spie),
    .io_dpath_status_upie(PTW_1_io_dpath_status_upie),
    .io_dpath_status_mie(PTW_1_io_dpath_status_mie),
    .io_dpath_status_hie(PTW_1_io_dpath_status_hie),
    .io_dpath_status_sie(PTW_1_io_dpath_status_sie),
    .io_dpath_status_uie(PTW_1_io_dpath_status_uie)
  );
  HellaCacheArbiter dcArb (
    .clk(dcArb_clk),
    .reset(dcArb_reset),
    .io_requestor_0_req_ready(dcArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_tag(dcArb_io_requestor_0_req_bits_tag),
    .io_requestor_0_req_bits_cmd(dcArb_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_typ(dcArb_io_requestor_0_req_bits_typ),
    .io_requestor_0_req_bits_phys(dcArb_io_requestor_0_req_bits_phys),
    .io_requestor_0_req_bits_data(dcArb_io_requestor_0_req_bits_data),
    .io_requestor_0_s1_kill(dcArb_io_requestor_0_s1_kill),
    .io_requestor_0_s1_data(dcArb_io_requestor_0_s1_data),
    .io_requestor_0_s2_nack(dcArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_addr(dcArb_io_requestor_0_resp_bits_addr),
    .io_requestor_0_resp_bits_tag(dcArb_io_requestor_0_resp_bits_tag),
    .io_requestor_0_resp_bits_cmd(dcArb_io_requestor_0_resp_bits_cmd),
    .io_requestor_0_resp_bits_typ(dcArb_io_requestor_0_resp_bits_typ),
    .io_requestor_0_resp_bits_data(dcArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_resp_bits_replay(dcArb_io_requestor_0_resp_bits_replay),
    .io_requestor_0_resp_bits_has_data(dcArb_io_requestor_0_resp_bits_has_data),
    .io_requestor_0_resp_bits_data_word_bypass(dcArb_io_requestor_0_resp_bits_data_word_bypass),
    .io_requestor_0_resp_bits_store_data(dcArb_io_requestor_0_resp_bits_store_data),
    .io_requestor_0_replay_next(dcArb_io_requestor_0_replay_next),
    .io_requestor_0_xcpt_ma_ld(dcArb_io_requestor_0_xcpt_ma_ld),
    .io_requestor_0_xcpt_ma_st(dcArb_io_requestor_0_xcpt_ma_st),
    .io_requestor_0_xcpt_pf_ld(dcArb_io_requestor_0_xcpt_pf_ld),
    .io_requestor_0_xcpt_pf_st(dcArb_io_requestor_0_xcpt_pf_st),
    .io_requestor_0_invalidate_lr(dcArb_io_requestor_0_invalidate_lr),
    .io_requestor_0_ordered(dcArb_io_requestor_0_ordered),
    .io_requestor_1_req_ready(dcArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_typ(dcArb_io_requestor_1_req_bits_typ),
    .io_requestor_1_req_bits_phys(dcArb_io_requestor_1_req_bits_phys),
    .io_requestor_1_req_bits_data(dcArb_io_requestor_1_req_bits_data),
    .io_requestor_1_s1_kill(dcArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data(dcArb_io_requestor_1_s1_data),
    .io_requestor_1_s2_nack(dcArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_addr(dcArb_io_requestor_1_resp_bits_addr),
    .io_requestor_1_resp_bits_tag(dcArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_cmd(dcArb_io_requestor_1_resp_bits_cmd),
    .io_requestor_1_resp_bits_typ(dcArb_io_requestor_1_resp_bits_typ),
    .io_requestor_1_resp_bits_data(dcArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_replay(dcArb_io_requestor_1_resp_bits_replay),
    .io_requestor_1_resp_bits_has_data(dcArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_resp_bits_data_word_bypass(dcArb_io_requestor_1_resp_bits_data_word_bypass),
    .io_requestor_1_resp_bits_store_data(dcArb_io_requestor_1_resp_bits_store_data),
    .io_requestor_1_replay_next(dcArb_io_requestor_1_replay_next),
    .io_requestor_1_xcpt_ma_ld(dcArb_io_requestor_1_xcpt_ma_ld),
    .io_requestor_1_xcpt_ma_st(dcArb_io_requestor_1_xcpt_ma_st),
    .io_requestor_1_xcpt_pf_ld(dcArb_io_requestor_1_xcpt_pf_ld),
    .io_requestor_1_xcpt_pf_st(dcArb_io_requestor_1_xcpt_pf_st),
    .io_requestor_1_invalidate_lr(dcArb_io_requestor_1_invalidate_lr),
    .io_requestor_1_ordered(dcArb_io_requestor_1_ordered),
    .io_mem_req_ready(dcArb_io_mem_req_ready),
    .io_mem_req_valid(dcArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcArb_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(dcArb_io_mem_req_bits_phys),
    .io_mem_req_bits_data(dcArb_io_mem_req_bits_data),
    .io_mem_s1_kill(dcArb_io_mem_s1_kill),
    .io_mem_s1_data(dcArb_io_mem_s1_data),
    .io_mem_s2_nack(dcArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcArb_io_mem_resp_valid),
    .io_mem_resp_bits_addr(dcArb_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(dcArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(dcArb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(dcArb_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(dcArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(dcArb_io_mem_resp_bits_store_data),
    .io_mem_replay_next(dcArb_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(dcArb_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(dcArb_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(dcArb_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(dcArb_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(dcArb_io_mem_invalidate_lr),
    .io_mem_ordered(dcArb_io_mem_ordered)
  );
  assign io_cached_0_acquire_valid = HellaCache_1_io_mem_acquire_valid;
  assign io_cached_0_acquire_bits_addr_block = HellaCache_1_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_bits_client_xact_id = HellaCache_1_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_beat = HellaCache_1_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_is_builtin_type = HellaCache_1_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_a_type = HellaCache_1_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_union = HellaCache_1_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_data = HellaCache_1_io_mem_acquire_bits_data;
  assign io_cached_0_probe_ready = HellaCache_1_io_mem_probe_ready;
  assign io_cached_0_release_valid = HellaCache_1_io_mem_release_valid;
  assign io_cached_0_release_bits_addr_beat = HellaCache_1_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_bits_addr_block = HellaCache_1_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_client_xact_id = HellaCache_1_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_voluntary = HellaCache_1_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_r_type = HellaCache_1_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_data = HellaCache_1_io_mem_release_bits_data;
  assign io_cached_0_grant_ready = HellaCache_1_io_mem_grant_ready;
  assign io_cached_0_finish_valid = HellaCache_1_io_mem_finish_valid;
  assign io_cached_0_finish_bits_manager_xact_id = HellaCache_1_io_mem_finish_bits_manager_xact_id;
  assign io_cached_0_finish_bits_manager_id = HellaCache_1_io_mem_finish_bits_manager_id;
  assign io_uncached_0_acquire_valid = uncachedArb_io_out_acquire_valid;
  assign io_uncached_0_acquire_bits_addr_block = uncachedArb_io_out_acquire_bits_addr_block;
  assign io_uncached_0_acquire_bits_client_xact_id = uncachedArb_io_out_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_beat = uncachedArb_io_out_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_is_builtin_type = uncachedArb_io_out_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_a_type = uncachedArb_io_out_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_union = uncachedArb_io_out_acquire_bits_union;
  assign io_uncached_0_acquire_bits_data = uncachedArb_io_out_acquire_bits_data;
  assign io_uncached_0_grant_ready = uncachedArb_io_out_grant_ready;
  assign core_clk = clk;
  assign core_reset = reset;
  assign core_io_prci_reset = io_prci_reset;
  assign core_io_prci_id = io_prci_id;
  assign core_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign core_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign core_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign core_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign core_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign core_io_imem_resp_valid = icache_io_cpu_resp_valid;
  assign core_io_imem_resp_bits_pc = icache_io_cpu_resp_bits_pc;
  assign core_io_imem_resp_bits_data_0 = icache_io_cpu_resp_bits_data_0;
  assign core_io_imem_resp_bits_mask = icache_io_cpu_resp_bits_mask;
  assign core_io_imem_resp_bits_xcpt_if = icache_io_cpu_resp_bits_xcpt_if;
  assign core_io_imem_btb_resp_valid = icache_io_cpu_btb_resp_valid;
  assign core_io_imem_btb_resp_bits_taken = icache_io_cpu_btb_resp_bits_taken;
  assign core_io_imem_btb_resp_bits_mask = icache_io_cpu_btb_resp_bits_mask;
  assign core_io_imem_btb_resp_bits_bridx = icache_io_cpu_btb_resp_bits_bridx;
  assign core_io_imem_btb_resp_bits_target = icache_io_cpu_btb_resp_bits_target;
  assign core_io_imem_btb_resp_bits_entry = icache_io_cpu_btb_resp_bits_entry;
  assign core_io_imem_btb_resp_bits_bht_history = icache_io_cpu_btb_resp_bits_bht_history;
  assign core_io_imem_btb_resp_bits_bht_value = icache_io_cpu_btb_resp_bits_bht_value;
  assign core_io_imem_npc = icache_io_cpu_npc;
  assign core_io_dmem_req_ready = dcArb_io_requestor_1_req_ready;
  assign core_io_dmem_s2_nack = dcArb_io_requestor_1_s2_nack;
  assign core_io_dmem_resp_valid = dcArb_io_requestor_1_resp_valid;
  assign core_io_dmem_resp_bits_addr = dcArb_io_requestor_1_resp_bits_addr;
  assign core_io_dmem_resp_bits_tag = dcArb_io_requestor_1_resp_bits_tag;
  assign core_io_dmem_resp_bits_cmd = dcArb_io_requestor_1_resp_bits_cmd;
  assign core_io_dmem_resp_bits_typ = dcArb_io_requestor_1_resp_bits_typ;
  assign core_io_dmem_resp_bits_data = dcArb_io_requestor_1_resp_bits_data;
  assign core_io_dmem_resp_bits_replay = dcArb_io_requestor_1_resp_bits_replay;
  assign core_io_dmem_resp_bits_has_data = dcArb_io_requestor_1_resp_bits_has_data;
  assign core_io_dmem_resp_bits_data_word_bypass = dcArb_io_requestor_1_resp_bits_data_word_bypass;
  assign core_io_dmem_resp_bits_store_data = dcArb_io_requestor_1_resp_bits_store_data;
  assign core_io_dmem_replay_next = dcArb_io_requestor_1_replay_next;
  assign core_io_dmem_xcpt_ma_ld = dcArb_io_requestor_1_xcpt_ma_ld;
  assign core_io_dmem_xcpt_ma_st = dcArb_io_requestor_1_xcpt_ma_st;
  assign core_io_dmem_xcpt_pf_ld = dcArb_io_requestor_1_xcpt_pf_ld;
  assign core_io_dmem_xcpt_pf_st = dcArb_io_requestor_1_xcpt_pf_st;
  assign core_io_dmem_ordered = dcArb_io_requestor_1_ordered;
  assign core_io_fpu_fcsr_flags_valid = GEN_0;
  assign core_io_fpu_fcsr_flags_bits = GEN_1;
  assign core_io_fpu_store_data = GEN_2;
  assign core_io_fpu_toint_data = GEN_3;
  assign core_io_fpu_fcsr_rdy = GEN_4;
  assign core_io_fpu_nack_mem = GEN_5;
  assign core_io_fpu_illegal_rm = GEN_6;
  assign core_io_fpu_dec_cmd = GEN_7;
  assign core_io_fpu_dec_ldst = GEN_8;
  assign core_io_fpu_dec_wen = GEN_9;
  assign core_io_fpu_dec_ren1 = GEN_10;
  assign core_io_fpu_dec_ren2 = GEN_11;
  assign core_io_fpu_dec_ren3 = GEN_12;
  assign core_io_fpu_dec_swap12 = GEN_13;
  assign core_io_fpu_dec_swap23 = GEN_14;
  assign core_io_fpu_dec_single = GEN_15;
  assign core_io_fpu_dec_fromint = GEN_16;
  assign core_io_fpu_dec_toint = GEN_17;
  assign core_io_fpu_dec_fastpipe = GEN_18;
  assign core_io_fpu_dec_fma = GEN_19;
  assign core_io_fpu_dec_div = GEN_20;
  assign core_io_fpu_dec_sqrt = GEN_21;
  assign core_io_fpu_dec_round = GEN_22;
  assign core_io_fpu_dec_wflags = GEN_23;
  assign core_io_fpu_sboard_set = GEN_24;
  assign core_io_fpu_sboard_clr = GEN_25;
  assign core_io_fpu_sboard_clra = GEN_26;
  assign core_io_fpu_cp_req_ready = GEN_27;
  assign core_io_fpu_cp_resp_valid = GEN_28;
  assign core_io_fpu_cp_resp_bits_data = GEN_29;
  assign core_io_fpu_cp_resp_bits_exc = GEN_30;
  assign core_io_rocc_cmd_ready = GEN_31;
  assign core_io_rocc_resp_valid = GEN_32;
  assign core_io_rocc_resp_bits_rd = GEN_33;
  assign core_io_rocc_resp_bits_data = GEN_34;
  assign core_io_rocc_mem_req_valid = GEN_35;
  assign core_io_rocc_mem_req_bits_addr = GEN_36;
  assign core_io_rocc_mem_req_bits_tag = GEN_37;
  assign core_io_rocc_mem_req_bits_cmd = GEN_38;
  assign core_io_rocc_mem_req_bits_typ = GEN_39;
  assign core_io_rocc_mem_req_bits_phys = GEN_40;
  assign core_io_rocc_mem_req_bits_data = GEN_41;
  assign core_io_rocc_mem_s1_kill = GEN_42;
  assign core_io_rocc_mem_s1_data = GEN_43;
  assign core_io_rocc_mem_invalidate_lr = GEN_44;
  assign core_io_rocc_busy = GEN_45;
  assign core_io_rocc_interrupt = GEN_46;
  assign core_io_rocc_autl_acquire_valid = GEN_47;
  assign core_io_rocc_autl_acquire_bits_addr_block = GEN_48;
  assign core_io_rocc_autl_acquire_bits_client_xact_id = GEN_49;
  assign core_io_rocc_autl_acquire_bits_addr_beat = GEN_50;
  assign core_io_rocc_autl_acquire_bits_is_builtin_type = GEN_51;
  assign core_io_rocc_autl_acquire_bits_a_type = GEN_52;
  assign core_io_rocc_autl_acquire_bits_union = GEN_53;
  assign core_io_rocc_autl_acquire_bits_data = GEN_54;
  assign core_io_rocc_autl_grant_ready = GEN_55;
  assign core_io_rocc_fpu_req_valid = GEN_56;
  assign core_io_rocc_fpu_req_bits_cmd = GEN_57;
  assign core_io_rocc_fpu_req_bits_ldst = GEN_58;
  assign core_io_rocc_fpu_req_bits_wen = GEN_59;
  assign core_io_rocc_fpu_req_bits_ren1 = GEN_60;
  assign core_io_rocc_fpu_req_bits_ren2 = GEN_61;
  assign core_io_rocc_fpu_req_bits_ren3 = GEN_62;
  assign core_io_rocc_fpu_req_bits_swap12 = GEN_63;
  assign core_io_rocc_fpu_req_bits_swap23 = GEN_64;
  assign core_io_rocc_fpu_req_bits_single = GEN_65;
  assign core_io_rocc_fpu_req_bits_fromint = GEN_66;
  assign core_io_rocc_fpu_req_bits_toint = GEN_67;
  assign core_io_rocc_fpu_req_bits_fastpipe = GEN_68;
  assign core_io_rocc_fpu_req_bits_fma = GEN_69;
  assign core_io_rocc_fpu_req_bits_div = GEN_70;
  assign core_io_rocc_fpu_req_bits_sqrt = GEN_71;
  assign core_io_rocc_fpu_req_bits_round = GEN_72;
  assign core_io_rocc_fpu_req_bits_wflags = GEN_73;
  assign core_io_rocc_fpu_req_bits_rm = GEN_74;
  assign core_io_rocc_fpu_req_bits_typ = GEN_75;
  assign core_io_rocc_fpu_req_bits_in1 = GEN_76;
  assign core_io_rocc_fpu_req_bits_in2 = GEN_77;
  assign core_io_rocc_fpu_req_bits_in3 = GEN_78;
  assign core_io_rocc_fpu_resp_ready = GEN_79;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_cpu_req_valid = core_io_imem_req_valid;
  assign icache_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
  assign icache_io_cpu_resp_ready = core_io_imem_resp_ready;
  assign icache_io_cpu_btb_update_valid = core_io_imem_btb_update_valid;
  assign icache_io_cpu_btb_update_bits_prediction_valid = core_io_imem_btb_update_bits_prediction_valid;
  assign icache_io_cpu_btb_update_bits_prediction_bits_taken = core_io_imem_btb_update_bits_prediction_bits_taken;
  assign icache_io_cpu_btb_update_bits_prediction_bits_mask = core_io_imem_btb_update_bits_prediction_bits_mask;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bridx = core_io_imem_btb_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_btb_update_bits_prediction_bits_target = core_io_imem_btb_update_bits_prediction_bits_target;
  assign icache_io_cpu_btb_update_bits_prediction_bits_entry = core_io_imem_btb_update_bits_prediction_bits_entry;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_history = core_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_value = core_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc;
  assign icache_io_cpu_btb_update_bits_target = core_io_imem_btb_update_bits_target;
  assign icache_io_cpu_btb_update_bits_taken = core_io_imem_btb_update_bits_taken;
  assign icache_io_cpu_btb_update_bits_isJump = core_io_imem_btb_update_bits_isJump;
  assign icache_io_cpu_btb_update_bits_isReturn = core_io_imem_btb_update_bits_isReturn;
  assign icache_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc;
  assign icache_io_cpu_bht_update_valid = core_io_imem_bht_update_valid;
  assign icache_io_cpu_bht_update_bits_prediction_valid = core_io_imem_bht_update_bits_prediction_valid;
  assign icache_io_cpu_bht_update_bits_prediction_bits_taken = core_io_imem_bht_update_bits_prediction_bits_taken;
  assign icache_io_cpu_bht_update_bits_prediction_bits_mask = core_io_imem_bht_update_bits_prediction_bits_mask;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bridx = core_io_imem_bht_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_bht_update_bits_prediction_bits_target = core_io_imem_bht_update_bits_prediction_bits_target;
  assign icache_io_cpu_bht_update_bits_prediction_bits_entry = core_io_imem_bht_update_bits_prediction_bits_entry;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_history = core_io_imem_bht_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_value = core_io_imem_bht_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc;
  assign icache_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken;
  assign icache_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict;
  assign icache_io_cpu_ras_update_valid = core_io_imem_ras_update_valid;
  assign icache_io_cpu_ras_update_bits_isCall = core_io_imem_ras_update_bits_isCall;
  assign icache_io_cpu_ras_update_bits_isReturn = core_io_imem_ras_update_bits_isReturn;
  assign icache_io_cpu_ras_update_bits_returnAddr = core_io_imem_ras_update_bits_returnAddr;
  assign icache_io_cpu_ras_update_bits_prediction_valid = core_io_imem_ras_update_bits_prediction_valid;
  assign icache_io_cpu_ras_update_bits_prediction_bits_taken = core_io_imem_ras_update_bits_prediction_bits_taken;
  assign icache_io_cpu_ras_update_bits_prediction_bits_mask = core_io_imem_ras_update_bits_prediction_bits_mask;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bridx = core_io_imem_ras_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_ras_update_bits_prediction_bits_target = core_io_imem_ras_update_bits_prediction_bits_target;
  assign icache_io_cpu_ras_update_bits_prediction_bits_entry = core_io_imem_ras_update_bits_prediction_bits_entry;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_history = core_io_imem_ras_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_value = core_io_imem_ras_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_flush_icache = core_io_imem_flush_icache;
  assign icache_io_cpu_flush_tlb = core_io_imem_flush_tlb;
  assign icache_io_ptw_req_ready = PTW_1_io_requestor_0_req_ready;
  assign icache_io_ptw_resp_valid = PTW_1_io_requestor_0_resp_valid;
  assign icache_io_ptw_resp_bits_pte_ppn = PTW_1_io_requestor_0_resp_bits_pte_ppn;
  assign icache_io_ptw_resp_bits_pte_reserved_for_software = PTW_1_io_requestor_0_resp_bits_pte_reserved_for_software;
  assign icache_io_ptw_resp_bits_pte_d = PTW_1_io_requestor_0_resp_bits_pte_d;
  assign icache_io_ptw_resp_bits_pte_r = PTW_1_io_requestor_0_resp_bits_pte_r;
  assign icache_io_ptw_resp_bits_pte_typ = PTW_1_io_requestor_0_resp_bits_pte_typ;
  assign icache_io_ptw_resp_bits_pte_v = PTW_1_io_requestor_0_resp_bits_pte_v;
  assign icache_io_ptw_ptbr_asid = PTW_1_io_requestor_0_ptbr_asid;
  assign icache_io_ptw_ptbr_ppn = PTW_1_io_requestor_0_ptbr_ppn;
  assign icache_io_ptw_invalidate = PTW_1_io_requestor_0_invalidate;
  assign icache_io_ptw_status_debug = PTW_1_io_requestor_0_status_debug;
  assign icache_io_ptw_status_prv = PTW_1_io_requestor_0_status_prv;
  assign icache_io_ptw_status_sd = PTW_1_io_requestor_0_status_sd;
  assign icache_io_ptw_status_zero3 = PTW_1_io_requestor_0_status_zero3;
  assign icache_io_ptw_status_sd_rv32 = PTW_1_io_requestor_0_status_sd_rv32;
  assign icache_io_ptw_status_zero2 = PTW_1_io_requestor_0_status_zero2;
  assign icache_io_ptw_status_vm = PTW_1_io_requestor_0_status_vm;
  assign icache_io_ptw_status_zero1 = PTW_1_io_requestor_0_status_zero1;
  assign icache_io_ptw_status_pum = PTW_1_io_requestor_0_status_pum;
  assign icache_io_ptw_status_mprv = PTW_1_io_requestor_0_status_mprv;
  assign icache_io_ptw_status_xs = PTW_1_io_requestor_0_status_xs;
  assign icache_io_ptw_status_fs = PTW_1_io_requestor_0_status_fs;
  assign icache_io_ptw_status_mpp = PTW_1_io_requestor_0_status_mpp;
  assign icache_io_ptw_status_hpp = PTW_1_io_requestor_0_status_hpp;
  assign icache_io_ptw_status_spp = PTW_1_io_requestor_0_status_spp;
  assign icache_io_ptw_status_mpie = PTW_1_io_requestor_0_status_mpie;
  assign icache_io_ptw_status_hpie = PTW_1_io_requestor_0_status_hpie;
  assign icache_io_ptw_status_spie = PTW_1_io_requestor_0_status_spie;
  assign icache_io_ptw_status_upie = PTW_1_io_requestor_0_status_upie;
  assign icache_io_ptw_status_mie = PTW_1_io_requestor_0_status_mie;
  assign icache_io_ptw_status_hie = PTW_1_io_requestor_0_status_hie;
  assign icache_io_ptw_status_sie = PTW_1_io_requestor_0_status_sie;
  assign icache_io_ptw_status_uie = PTW_1_io_requestor_0_status_uie;
  assign icache_io_mem_acquire_ready = uncachedArb_io_in_0_acquire_ready;
  assign icache_io_mem_grant_valid = uncachedArb_io_in_0_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = uncachedArb_io_in_0_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = uncachedArb_io_in_0_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = uncachedArb_io_in_0_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = uncachedArb_io_in_0_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = uncachedArb_io_in_0_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = uncachedArb_io_in_0_grant_bits_data;
  assign HellaCache_1_clk = clk;
  assign HellaCache_1_reset = reset;
  assign HellaCache_1_io_cpu_req_valid = dcArb_io_mem_req_valid;
  assign HellaCache_1_io_cpu_req_bits_addr = dcArb_io_mem_req_bits_addr;
  assign HellaCache_1_io_cpu_req_bits_tag = dcArb_io_mem_req_bits_tag;
  assign HellaCache_1_io_cpu_req_bits_cmd = dcArb_io_mem_req_bits_cmd;
  assign HellaCache_1_io_cpu_req_bits_typ = dcArb_io_mem_req_bits_typ;
  assign HellaCache_1_io_cpu_req_bits_phys = dcArb_io_mem_req_bits_phys;
  assign HellaCache_1_io_cpu_req_bits_data = dcArb_io_mem_req_bits_data;
  assign HellaCache_1_io_cpu_s1_kill = dcArb_io_mem_s1_kill;
  assign HellaCache_1_io_cpu_s1_data = dcArb_io_mem_s1_data;
  assign HellaCache_1_io_cpu_invalidate_lr = dcArb_io_mem_invalidate_lr;
  assign HellaCache_1_io_ptw_req_ready = PTW_1_io_requestor_1_req_ready;
  assign HellaCache_1_io_ptw_resp_valid = PTW_1_io_requestor_1_resp_valid;
  assign HellaCache_1_io_ptw_resp_bits_pte_ppn = PTW_1_io_requestor_1_resp_bits_pte_ppn;
  assign HellaCache_1_io_ptw_resp_bits_pte_reserved_for_software = PTW_1_io_requestor_1_resp_bits_pte_reserved_for_software;
  assign HellaCache_1_io_ptw_resp_bits_pte_d = PTW_1_io_requestor_1_resp_bits_pte_d;
  assign HellaCache_1_io_ptw_resp_bits_pte_r = PTW_1_io_requestor_1_resp_bits_pte_r;
  assign HellaCache_1_io_ptw_resp_bits_pte_typ = PTW_1_io_requestor_1_resp_bits_pte_typ;
  assign HellaCache_1_io_ptw_resp_bits_pte_v = PTW_1_io_requestor_1_resp_bits_pte_v;
  assign HellaCache_1_io_ptw_ptbr_asid = PTW_1_io_requestor_1_ptbr_asid;
  assign HellaCache_1_io_ptw_ptbr_ppn = PTW_1_io_requestor_1_ptbr_ppn;
  assign HellaCache_1_io_ptw_invalidate = PTW_1_io_requestor_1_invalidate;
  assign HellaCache_1_io_ptw_status_debug = PTW_1_io_requestor_1_status_debug;
  assign HellaCache_1_io_ptw_status_prv = PTW_1_io_requestor_1_status_prv;
  assign HellaCache_1_io_ptw_status_sd = PTW_1_io_requestor_1_status_sd;
  assign HellaCache_1_io_ptw_status_zero3 = PTW_1_io_requestor_1_status_zero3;
  assign HellaCache_1_io_ptw_status_sd_rv32 = PTW_1_io_requestor_1_status_sd_rv32;
  assign HellaCache_1_io_ptw_status_zero2 = PTW_1_io_requestor_1_status_zero2;
  assign HellaCache_1_io_ptw_status_vm = PTW_1_io_requestor_1_status_vm;
  assign HellaCache_1_io_ptw_status_zero1 = PTW_1_io_requestor_1_status_zero1;
  assign HellaCache_1_io_ptw_status_pum = PTW_1_io_requestor_1_status_pum;
  assign HellaCache_1_io_ptw_status_mprv = PTW_1_io_requestor_1_status_mprv;
  assign HellaCache_1_io_ptw_status_xs = PTW_1_io_requestor_1_status_xs;
  assign HellaCache_1_io_ptw_status_fs = PTW_1_io_requestor_1_status_fs;
  assign HellaCache_1_io_ptw_status_mpp = PTW_1_io_requestor_1_status_mpp;
  assign HellaCache_1_io_ptw_status_hpp = PTW_1_io_requestor_1_status_hpp;
  assign HellaCache_1_io_ptw_status_spp = PTW_1_io_requestor_1_status_spp;
  assign HellaCache_1_io_ptw_status_mpie = PTW_1_io_requestor_1_status_mpie;
  assign HellaCache_1_io_ptw_status_hpie = PTW_1_io_requestor_1_status_hpie;
  assign HellaCache_1_io_ptw_status_spie = PTW_1_io_requestor_1_status_spie;
  assign HellaCache_1_io_ptw_status_upie = PTW_1_io_requestor_1_status_upie;
  assign HellaCache_1_io_ptw_status_mie = PTW_1_io_requestor_1_status_mie;
  assign HellaCache_1_io_ptw_status_hie = PTW_1_io_requestor_1_status_hie;
  assign HellaCache_1_io_ptw_status_sie = PTW_1_io_requestor_1_status_sie;
  assign HellaCache_1_io_ptw_status_uie = PTW_1_io_requestor_1_status_uie;
  assign HellaCache_1_io_mem_acquire_ready = io_cached_0_acquire_ready;
  assign HellaCache_1_io_mem_probe_valid = io_cached_0_probe_valid;
  assign HellaCache_1_io_mem_probe_bits_addr_block = io_cached_0_probe_bits_addr_block;
  assign HellaCache_1_io_mem_probe_bits_p_type = io_cached_0_probe_bits_p_type;
  assign HellaCache_1_io_mem_release_ready = io_cached_0_release_ready;
  assign HellaCache_1_io_mem_grant_valid = io_cached_0_grant_valid;
  assign HellaCache_1_io_mem_grant_bits_addr_beat = io_cached_0_grant_bits_addr_beat;
  assign HellaCache_1_io_mem_grant_bits_client_xact_id = io_cached_0_grant_bits_client_xact_id;
  assign HellaCache_1_io_mem_grant_bits_manager_xact_id = io_cached_0_grant_bits_manager_xact_id;
  assign HellaCache_1_io_mem_grant_bits_is_builtin_type = io_cached_0_grant_bits_is_builtin_type;
  assign HellaCache_1_io_mem_grant_bits_g_type = io_cached_0_grant_bits_g_type;
  assign HellaCache_1_io_mem_grant_bits_data = io_cached_0_grant_bits_data;
  assign HellaCache_1_io_mem_grant_bits_manager_id = io_cached_0_grant_bits_manager_id;
  assign HellaCache_1_io_mem_finish_ready = io_cached_0_finish_ready;
  assign uncachedArb_clk = clk;
  assign uncachedArb_reset = reset;
  assign uncachedArb_io_in_0_acquire_valid = icache_io_mem_acquire_valid;
  assign uncachedArb_io_in_0_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign uncachedArb_io_in_0_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign uncachedArb_io_in_0_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign uncachedArb_io_in_0_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign uncachedArb_io_in_0_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign uncachedArb_io_in_0_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign uncachedArb_io_in_0_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign uncachedArb_io_in_0_grant_ready = icache_io_mem_grant_ready;
  assign uncachedArb_io_out_acquire_ready = io_uncached_0_acquire_ready;
  assign uncachedArb_io_out_grant_valid = io_uncached_0_grant_valid;
  assign uncachedArb_io_out_grant_bits_addr_beat = io_uncached_0_grant_bits_addr_beat;
  assign uncachedArb_io_out_grant_bits_client_xact_id = io_uncached_0_grant_bits_client_xact_id;
  assign uncachedArb_io_out_grant_bits_manager_xact_id = io_uncached_0_grant_bits_manager_xact_id;
  assign uncachedArb_io_out_grant_bits_is_builtin_type = io_uncached_0_grant_bits_is_builtin_type;
  assign uncachedArb_io_out_grant_bits_g_type = io_uncached_0_grant_bits_g_type;
  assign uncachedArb_io_out_grant_bits_data = io_uncached_0_grant_bits_data;
  assign PTW_1_clk = clk;
  assign PTW_1_reset = reset;
  assign PTW_1_io_requestor_0_req_valid = icache_io_ptw_req_valid;
  assign PTW_1_io_requestor_0_req_bits_addr = icache_io_ptw_req_bits_addr;
  assign PTW_1_io_requestor_0_req_bits_prv = icache_io_ptw_req_bits_prv;
  assign PTW_1_io_requestor_0_req_bits_store = icache_io_ptw_req_bits_store;
  assign PTW_1_io_requestor_0_req_bits_fetch = icache_io_ptw_req_bits_fetch;
  assign PTW_1_io_requestor_1_req_valid = HellaCache_1_io_ptw_req_valid;
  assign PTW_1_io_requestor_1_req_bits_addr = HellaCache_1_io_ptw_req_bits_addr;
  assign PTW_1_io_requestor_1_req_bits_prv = HellaCache_1_io_ptw_req_bits_prv;
  assign PTW_1_io_requestor_1_req_bits_store = HellaCache_1_io_ptw_req_bits_store;
  assign PTW_1_io_requestor_1_req_bits_fetch = HellaCache_1_io_ptw_req_bits_fetch;
  assign PTW_1_io_mem_req_ready = dcArb_io_requestor_0_req_ready;
  assign PTW_1_io_mem_s2_nack = dcArb_io_requestor_0_s2_nack;
  assign PTW_1_io_mem_resp_valid = dcArb_io_requestor_0_resp_valid;
  assign PTW_1_io_mem_resp_bits_addr = dcArb_io_requestor_0_resp_bits_addr;
  assign PTW_1_io_mem_resp_bits_tag = dcArb_io_requestor_0_resp_bits_tag;
  assign PTW_1_io_mem_resp_bits_cmd = dcArb_io_requestor_0_resp_bits_cmd;
  assign PTW_1_io_mem_resp_bits_typ = dcArb_io_requestor_0_resp_bits_typ;
  assign PTW_1_io_mem_resp_bits_data = dcArb_io_requestor_0_resp_bits_data;
  assign PTW_1_io_mem_resp_bits_replay = dcArb_io_requestor_0_resp_bits_replay;
  assign PTW_1_io_mem_resp_bits_has_data = dcArb_io_requestor_0_resp_bits_has_data;
  assign PTW_1_io_mem_resp_bits_data_word_bypass = dcArb_io_requestor_0_resp_bits_data_word_bypass;
  assign PTW_1_io_mem_resp_bits_store_data = dcArb_io_requestor_0_resp_bits_store_data;
  assign PTW_1_io_mem_replay_next = dcArb_io_requestor_0_replay_next;
  assign PTW_1_io_mem_xcpt_ma_ld = dcArb_io_requestor_0_xcpt_ma_ld;
  assign PTW_1_io_mem_xcpt_ma_st = dcArb_io_requestor_0_xcpt_ma_st;
  assign PTW_1_io_mem_xcpt_pf_ld = dcArb_io_requestor_0_xcpt_pf_ld;
  assign PTW_1_io_mem_xcpt_pf_st = dcArb_io_requestor_0_xcpt_pf_st;
  assign PTW_1_io_mem_ordered = dcArb_io_requestor_0_ordered;
  assign PTW_1_io_dpath_ptbr_asid = core_io_ptw_ptbr_asid;
  assign PTW_1_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn;
  assign PTW_1_io_dpath_invalidate = core_io_ptw_invalidate;
  assign PTW_1_io_dpath_status_debug = core_io_ptw_status_debug;
  assign PTW_1_io_dpath_status_prv = core_io_ptw_status_prv;
  assign PTW_1_io_dpath_status_sd = core_io_ptw_status_sd;
  assign PTW_1_io_dpath_status_zero3 = core_io_ptw_status_zero3;
  assign PTW_1_io_dpath_status_sd_rv32 = core_io_ptw_status_sd_rv32;
  assign PTW_1_io_dpath_status_zero2 = core_io_ptw_status_zero2;
  assign PTW_1_io_dpath_status_vm = core_io_ptw_status_vm;
  assign PTW_1_io_dpath_status_zero1 = core_io_ptw_status_zero1;
  assign PTW_1_io_dpath_status_pum = core_io_ptw_status_pum;
  assign PTW_1_io_dpath_status_mprv = core_io_ptw_status_mprv;
  assign PTW_1_io_dpath_status_xs = core_io_ptw_status_xs;
  assign PTW_1_io_dpath_status_fs = core_io_ptw_status_fs;
  assign PTW_1_io_dpath_status_mpp = core_io_ptw_status_mpp;
  assign PTW_1_io_dpath_status_hpp = core_io_ptw_status_hpp;
  assign PTW_1_io_dpath_status_spp = core_io_ptw_status_spp;
  assign PTW_1_io_dpath_status_mpie = core_io_ptw_status_mpie;
  assign PTW_1_io_dpath_status_hpie = core_io_ptw_status_hpie;
  assign PTW_1_io_dpath_status_spie = core_io_ptw_status_spie;
  assign PTW_1_io_dpath_status_upie = core_io_ptw_status_upie;
  assign PTW_1_io_dpath_status_mie = core_io_ptw_status_mie;
  assign PTW_1_io_dpath_status_hie = core_io_ptw_status_hie;
  assign PTW_1_io_dpath_status_sie = core_io_ptw_status_sie;
  assign PTW_1_io_dpath_status_uie = core_io_ptw_status_uie;
  assign dcArb_clk = clk;
  assign dcArb_reset = reset;
  assign dcArb_io_requestor_0_req_valid = PTW_1_io_mem_req_valid;
  assign dcArb_io_requestor_0_req_bits_addr = PTW_1_io_mem_req_bits_addr;
  assign dcArb_io_requestor_0_req_bits_tag = PTW_1_io_mem_req_bits_tag;
  assign dcArb_io_requestor_0_req_bits_cmd = PTW_1_io_mem_req_bits_cmd;
  assign dcArb_io_requestor_0_req_bits_typ = PTW_1_io_mem_req_bits_typ;
  assign dcArb_io_requestor_0_req_bits_phys = PTW_1_io_mem_req_bits_phys;
  assign dcArb_io_requestor_0_req_bits_data = PTW_1_io_mem_req_bits_data;
  assign dcArb_io_requestor_0_s1_kill = PTW_1_io_mem_s1_kill;
  assign dcArb_io_requestor_0_s1_data = PTW_1_io_mem_s1_data;
  assign dcArb_io_requestor_0_invalidate_lr = PTW_1_io_mem_invalidate_lr;
  assign dcArb_io_requestor_1_req_valid = core_io_dmem_req_valid;
  assign dcArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr;
  assign dcArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag;
  assign dcArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd;
  assign dcArb_io_requestor_1_req_bits_typ = core_io_dmem_req_bits_typ;
  assign dcArb_io_requestor_1_req_bits_phys = core_io_dmem_req_bits_phys;
  assign dcArb_io_requestor_1_req_bits_data = core_io_dmem_req_bits_data;
  assign dcArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill;
  assign dcArb_io_requestor_1_s1_data = core_io_dmem_s1_data;
  assign dcArb_io_requestor_1_invalidate_lr = core_io_dmem_invalidate_lr;
  assign dcArb_io_mem_req_ready = HellaCache_1_io_cpu_req_ready;
  assign dcArb_io_mem_s2_nack = HellaCache_1_io_cpu_s2_nack;
  assign dcArb_io_mem_resp_valid = HellaCache_1_io_cpu_resp_valid;
  assign dcArb_io_mem_resp_bits_addr = HellaCache_1_io_cpu_resp_bits_addr;
  assign dcArb_io_mem_resp_bits_tag = HellaCache_1_io_cpu_resp_bits_tag;
  assign dcArb_io_mem_resp_bits_cmd = HellaCache_1_io_cpu_resp_bits_cmd;
  assign dcArb_io_mem_resp_bits_typ = HellaCache_1_io_cpu_resp_bits_typ;
  assign dcArb_io_mem_resp_bits_data = HellaCache_1_io_cpu_resp_bits_data;
  assign dcArb_io_mem_resp_bits_replay = HellaCache_1_io_cpu_resp_bits_replay;
  assign dcArb_io_mem_resp_bits_has_data = HellaCache_1_io_cpu_resp_bits_has_data;
  assign dcArb_io_mem_resp_bits_data_word_bypass = HellaCache_1_io_cpu_resp_bits_data_word_bypass;
  assign dcArb_io_mem_resp_bits_store_data = HellaCache_1_io_cpu_resp_bits_store_data;
  assign dcArb_io_mem_replay_next = HellaCache_1_io_cpu_replay_next;
  assign dcArb_io_mem_xcpt_ma_ld = HellaCache_1_io_cpu_xcpt_ma_ld;
  assign dcArb_io_mem_xcpt_ma_st = HellaCache_1_io_cpu_xcpt_ma_st;
  assign dcArb_io_mem_xcpt_pf_ld = HellaCache_1_io_cpu_xcpt_pf_ld;
  assign dcArb_io_mem_xcpt_pf_st = HellaCache_1_io_cpu_xcpt_pf_st;
  assign dcArb_io_mem_ordered = HellaCache_1_io_cpu_ordered;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_80 = {1{$random}};
  GEN_0 = GEN_80[0:0];
  GEN_81 = {1{$random}};
  GEN_1 = GEN_81[4:0];
  GEN_82 = {2{$random}};
  GEN_2 = GEN_82[63:0];
  GEN_83 = {2{$random}};
  GEN_3 = GEN_83[63:0];
  GEN_84 = {1{$random}};
  GEN_4 = GEN_84[0:0];
  GEN_85 = {1{$random}};
  GEN_5 = GEN_85[0:0];
  GEN_86 = {1{$random}};
  GEN_6 = GEN_86[0:0];
  GEN_87 = {1{$random}};
  GEN_7 = GEN_87[4:0];
  GEN_88 = {1{$random}};
  GEN_8 = GEN_88[0:0];
  GEN_89 = {1{$random}};
  GEN_9 = GEN_89[0:0];
  GEN_90 = {1{$random}};
  GEN_10 = GEN_90[0:0];
  GEN_91 = {1{$random}};
  GEN_11 = GEN_91[0:0];
  GEN_92 = {1{$random}};
  GEN_12 = GEN_92[0:0];
  GEN_93 = {1{$random}};
  GEN_13 = GEN_93[0:0];
  GEN_94 = {1{$random}};
  GEN_14 = GEN_94[0:0];
  GEN_95 = {1{$random}};
  GEN_15 = GEN_95[0:0];
  GEN_96 = {1{$random}};
  GEN_16 = GEN_96[0:0];
  GEN_97 = {1{$random}};
  GEN_17 = GEN_97[0:0];
  GEN_98 = {1{$random}};
  GEN_18 = GEN_98[0:0];
  GEN_99 = {1{$random}};
  GEN_19 = GEN_99[0:0];
  GEN_100 = {1{$random}};
  GEN_20 = GEN_100[0:0];
  GEN_101 = {1{$random}};
  GEN_21 = GEN_101[0:0];
  GEN_102 = {1{$random}};
  GEN_22 = GEN_102[0:0];
  GEN_103 = {1{$random}};
  GEN_23 = GEN_103[0:0];
  GEN_104 = {1{$random}};
  GEN_24 = GEN_104[0:0];
  GEN_105 = {1{$random}};
  GEN_25 = GEN_105[0:0];
  GEN_106 = {1{$random}};
  GEN_26 = GEN_106[4:0];
  GEN_107 = {1{$random}};
  GEN_27 = GEN_107[0:0];
  GEN_108 = {1{$random}};
  GEN_28 = GEN_108[0:0];
  GEN_109 = {3{$random}};
  GEN_29 = GEN_109[64:0];
  GEN_110 = {1{$random}};
  GEN_30 = GEN_110[4:0];
  GEN_111 = {1{$random}};
  GEN_31 = GEN_111[0:0];
  GEN_112 = {1{$random}};
  GEN_32 = GEN_112[0:0];
  GEN_113 = {1{$random}};
  GEN_33 = GEN_113[4:0];
  GEN_114 = {2{$random}};
  GEN_34 = GEN_114[63:0];
  GEN_115 = {1{$random}};
  GEN_35 = GEN_115[0:0];
  GEN_116 = {2{$random}};
  GEN_36 = GEN_116[39:0];
  GEN_117 = {1{$random}};
  GEN_37 = GEN_117[8:0];
  GEN_118 = {1{$random}};
  GEN_38 = GEN_118[4:0];
  GEN_119 = {1{$random}};
  GEN_39 = GEN_119[2:0];
  GEN_120 = {1{$random}};
  GEN_40 = GEN_120[0:0];
  GEN_121 = {2{$random}};
  GEN_41 = GEN_121[63:0];
  GEN_122 = {1{$random}};
  GEN_42 = GEN_122[0:0];
  GEN_123 = {2{$random}};
  GEN_43 = GEN_123[63:0];
  GEN_124 = {1{$random}};
  GEN_44 = GEN_124[0:0];
  GEN_125 = {1{$random}};
  GEN_45 = GEN_125[0:0];
  GEN_126 = {1{$random}};
  GEN_46 = GEN_126[0:0];
  GEN_127 = {1{$random}};
  GEN_47 = GEN_127[0:0];
  GEN_128 = {1{$random}};
  GEN_48 = GEN_128[25:0];
  GEN_129 = {1{$random}};
  GEN_49 = GEN_129[1:0];
  GEN_130 = {1{$random}};
  GEN_50 = GEN_130[2:0];
  GEN_131 = {1{$random}};
  GEN_51 = GEN_131[0:0];
  GEN_132 = {1{$random}};
  GEN_52 = GEN_132[2:0];
  GEN_133 = {1{$random}};
  GEN_53 = GEN_133[11:0];
  GEN_134 = {2{$random}};
  GEN_54 = GEN_134[63:0];
  GEN_135 = {1{$random}};
  GEN_55 = GEN_135[0:0];
  GEN_136 = {1{$random}};
  GEN_56 = GEN_136[0:0];
  GEN_137 = {1{$random}};
  GEN_57 = GEN_137[4:0];
  GEN_138 = {1{$random}};
  GEN_58 = GEN_138[0:0];
  GEN_139 = {1{$random}};
  GEN_59 = GEN_139[0:0];
  GEN_140 = {1{$random}};
  GEN_60 = GEN_140[0:0];
  GEN_141 = {1{$random}};
  GEN_61 = GEN_141[0:0];
  GEN_142 = {1{$random}};
  GEN_62 = GEN_142[0:0];
  GEN_143 = {1{$random}};
  GEN_63 = GEN_143[0:0];
  GEN_144 = {1{$random}};
  GEN_64 = GEN_144[0:0];
  GEN_145 = {1{$random}};
  GEN_65 = GEN_145[0:0];
  GEN_146 = {1{$random}};
  GEN_66 = GEN_146[0:0];
  GEN_147 = {1{$random}};
  GEN_67 = GEN_147[0:0];
  GEN_148 = {1{$random}};
  GEN_68 = GEN_148[0:0];
  GEN_149 = {1{$random}};
  GEN_69 = GEN_149[0:0];
  GEN_150 = {1{$random}};
  GEN_70 = GEN_150[0:0];
  GEN_151 = {1{$random}};
  GEN_71 = GEN_151[0:0];
  GEN_152 = {1{$random}};
  GEN_72 = GEN_152[0:0];
  GEN_153 = {1{$random}};
  GEN_73 = GEN_153[0:0];
  GEN_154 = {1{$random}};
  GEN_74 = GEN_154[2:0];
  GEN_155 = {1{$random}};
  GEN_75 = GEN_155[1:0];
  GEN_156 = {3{$random}};
  GEN_76 = GEN_156[64:0];
  GEN_157 = {3{$random}};
  GEN_77 = GEN_157[64:0];
  GEN_158 = {3{$random}};
  GEN_78 = GEN_158[64:0];
  GEN_159 = {1{$random}};
  GEN_79 = GEN_159[0:0];
  end
`endif
endmodule
module Queue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input   io_enq_bits_payload_is_builtin_type,
  input  [2:0] io_enq_bits_payload_a_type,
  input  [11:0] io_enq_bits_payload_union,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output [2:0] io_deq_bits_payload_addr_beat,
  output  io_deq_bits_payload_is_builtin_type,
  output [2:0] io_deq_bits_payload_a_type,
  output [11:0] io_deq_bits_payload_union,
  output [63:0] io_deq_bits_payload_data,
  output  io_count
);
  reg [1:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1294_data;
  wire  ram_header_src_T_1294_addr;
  wire  ram_header_src_T_1294_en;
  wire [1:0] ram_header_src_T_1160_data;
  wire  ram_header_src_T_1160_addr;
  wire  ram_header_src_T_1160_mask;
  wire  ram_header_src_T_1160_en;
  reg [1:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1294_data;
  wire  ram_header_dst_T_1294_addr;
  wire  ram_header_dst_T_1294_en;
  wire [1:0] ram_header_dst_T_1160_data;
  wire  ram_header_dst_T_1160_addr;
  wire  ram_header_dst_T_1160_mask;
  wire  ram_header_dst_T_1160_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1294_data;
  wire  ram_payload_addr_block_T_1294_addr;
  wire  ram_payload_addr_block_T_1294_en;
  wire [25:0] ram_payload_addr_block_T_1160_data;
  wire  ram_payload_addr_block_T_1160_addr;
  wire  ram_payload_addr_block_T_1160_mask;
  wire  ram_payload_addr_block_T_1160_en;
  reg [1:0] ram_payload_client_xact_id [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_client_xact_id_T_1294_data;
  wire  ram_payload_client_xact_id_T_1294_addr;
  wire  ram_payload_client_xact_id_T_1294_en;
  wire [1:0] ram_payload_client_xact_id_T_1160_data;
  wire  ram_payload_client_xact_id_T_1160_addr;
  wire  ram_payload_client_xact_id_T_1160_mask;
  wire  ram_payload_client_xact_id_T_1160_en;
  reg [2:0] ram_payload_addr_beat [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_payload_addr_beat_T_1294_data;
  wire  ram_payload_addr_beat_T_1294_addr;
  wire  ram_payload_addr_beat_T_1294_en;
  wire [2:0] ram_payload_addr_beat_T_1160_data;
  wire  ram_payload_addr_beat_T_1160_addr;
  wire  ram_payload_addr_beat_T_1160_mask;
  wire  ram_payload_addr_beat_T_1160_en;
  reg  ram_payload_is_builtin_type [0:0];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1294_data;
  wire  ram_payload_is_builtin_type_T_1294_addr;
  wire  ram_payload_is_builtin_type_T_1294_en;
  wire  ram_payload_is_builtin_type_T_1160_data;
  wire  ram_payload_is_builtin_type_T_1160_addr;
  wire  ram_payload_is_builtin_type_T_1160_mask;
  wire  ram_payload_is_builtin_type_T_1160_en;
  reg [2:0] ram_payload_a_type [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_a_type_T_1294_data;
  wire  ram_payload_a_type_T_1294_addr;
  wire  ram_payload_a_type_T_1294_en;
  wire [2:0] ram_payload_a_type_T_1160_data;
  wire  ram_payload_a_type_T_1160_addr;
  wire  ram_payload_a_type_T_1160_mask;
  wire  ram_payload_a_type_T_1160_en;
  reg [11:0] ram_payload_union [0:0];
  reg [31:0] GEN_7;
  wire [11:0] ram_payload_union_T_1294_data;
  wire  ram_payload_union_T_1294_addr;
  wire  ram_payload_union_T_1294_en;
  wire [11:0] ram_payload_union_T_1160_data;
  wire  ram_payload_union_T_1160_addr;
  wire  ram_payload_union_T_1160_mask;
  wire  ram_payload_union_T_1160_en;
  reg [63:0] ram_payload_data [0:0];
  reg [63:0] GEN_8;
  wire [63:0] ram_payload_data_T_1294_data;
  wire  ram_payload_data_T_1294_addr;
  wire  ram_payload_data_T_1294_en;
  wire [63:0] ram_payload_data_T_1160_data;
  wire  ram_payload_data_T_1160_addr;
  wire  ram_payload_data_T_1160_mask;
  wire  ram_payload_data_T_1160_en;
  reg  maybe_full;
  reg [31:0] GEN_9;
  wire  T_1157;
  wire  T_1158;
  wire  do_enq;
  wire  T_1159;
  wire  do_deq;
  wire  T_1289;
  wire  GEN_21;
  wire  T_1291;
  wire [1:0] T_1421;
  wire  ptr_diff;
  wire [1:0] T_1423;
  assign io_enq_ready = T_1157;
  assign io_deq_valid = T_1291;
  assign io_deq_bits_header_src = ram_header_src_T_1294_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1294_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1294_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1294_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1294_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1294_data;
  assign io_deq_bits_payload_a_type = ram_payload_a_type_T_1294_data;
  assign io_deq_bits_payload_union = ram_payload_union_T_1294_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1294_data;
  assign io_count = T_1423[0];
  assign ram_header_src_T_1294_addr = 1'h0;
  assign ram_header_src_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_src_T_1294_data = ram_header_src[ram_header_src_T_1294_addr];
  `else
  assign ram_header_src_T_1294_data = ram_header_src_T_1294_addr >= 1'h1 ? $random : ram_header_src[ram_header_src_T_1294_addr];
  `endif
  assign ram_header_src_T_1160_data = io_enq_bits_header_src;
  assign ram_header_src_T_1160_addr = 1'h0;
  assign ram_header_src_T_1160_mask = do_enq;
  assign ram_header_src_T_1160_en = do_enq;
  assign ram_header_dst_T_1294_addr = 1'h0;
  assign ram_header_dst_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_dst_T_1294_data = ram_header_dst[ram_header_dst_T_1294_addr];
  `else
  assign ram_header_dst_T_1294_data = ram_header_dst_T_1294_addr >= 1'h1 ? $random : ram_header_dst[ram_header_dst_T_1294_addr];
  `endif
  assign ram_header_dst_T_1160_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1160_addr = 1'h0;
  assign ram_header_dst_T_1160_mask = do_enq;
  assign ram_header_dst_T_1160_en = do_enq;
  assign ram_payload_addr_block_T_1294_addr = 1'h0;
  assign ram_payload_addr_block_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_block_T_1294_data = ram_payload_addr_block[ram_payload_addr_block_T_1294_addr];
  `else
  assign ram_payload_addr_block_T_1294_data = ram_payload_addr_block_T_1294_addr >= 1'h1 ? $random : ram_payload_addr_block[ram_payload_addr_block_T_1294_addr];
  `endif
  assign ram_payload_addr_block_T_1160_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1160_addr = 1'h0;
  assign ram_payload_addr_block_T_1160_mask = do_enq;
  assign ram_payload_addr_block_T_1160_en = do_enq;
  assign ram_payload_client_xact_id_T_1294_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `else
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id_T_1294_addr >= 1'h1 ? $random : ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `endif
  assign ram_payload_client_xact_id_T_1160_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1160_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1160_mask = do_enq;
  assign ram_payload_client_xact_id_T_1160_en = do_enq;
  assign ram_payload_addr_beat_T_1294_addr = 1'h0;
  assign ram_payload_addr_beat_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `else
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat_T_1294_addr >= 1'h1 ? $random : ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `endif
  assign ram_payload_addr_beat_T_1160_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1160_addr = 1'h0;
  assign ram_payload_addr_beat_T_1160_mask = do_enq;
  assign ram_payload_addr_beat_T_1160_en = do_enq;
  assign ram_payload_is_builtin_type_T_1294_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_is_builtin_type_T_1294_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1294_addr];
  `else
  assign ram_payload_is_builtin_type_T_1294_data = ram_payload_is_builtin_type_T_1294_addr >= 1'h1 ? $random : ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1294_addr];
  `endif
  assign ram_payload_is_builtin_type_T_1160_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1160_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1160_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1160_en = do_enq;
  assign ram_payload_a_type_T_1294_addr = 1'h0;
  assign ram_payload_a_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_a_type_T_1294_data = ram_payload_a_type[ram_payload_a_type_T_1294_addr];
  `else
  assign ram_payload_a_type_T_1294_data = ram_payload_a_type_T_1294_addr >= 1'h1 ? $random : ram_payload_a_type[ram_payload_a_type_T_1294_addr];
  `endif
  assign ram_payload_a_type_T_1160_data = io_enq_bits_payload_a_type;
  assign ram_payload_a_type_T_1160_addr = 1'h0;
  assign ram_payload_a_type_T_1160_mask = do_enq;
  assign ram_payload_a_type_T_1160_en = do_enq;
  assign ram_payload_union_T_1294_addr = 1'h0;
  assign ram_payload_union_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_union_T_1294_data = ram_payload_union[ram_payload_union_T_1294_addr];
  `else
  assign ram_payload_union_T_1294_data = ram_payload_union_T_1294_addr >= 1'h1 ? $random : ram_payload_union[ram_payload_union_T_1294_addr];
  `endif
  assign ram_payload_union_T_1160_data = io_enq_bits_payload_union;
  assign ram_payload_union_T_1160_addr = 1'h0;
  assign ram_payload_union_T_1160_mask = do_enq;
  assign ram_payload_union_T_1160_en = do_enq;
  assign ram_payload_data_T_1294_addr = 1'h0;
  assign ram_payload_data_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_data_T_1294_data = ram_payload_data[ram_payload_data_T_1294_addr];
  `else
  assign ram_payload_data_T_1294_data = ram_payload_data_T_1294_addr >= 1'h1 ? $random : ram_payload_data[ram_payload_data_T_1294_addr];
  `endif
  assign ram_payload_data_T_1160_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1160_addr = 1'h0;
  assign ram_payload_data_T_1160_mask = do_enq;
  assign ram_payload_data_T_1160_en = do_enq;
  assign T_1157 = maybe_full == 1'h0;
  assign T_1158 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1158;
  assign T_1159 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1159;
  assign T_1289 = do_enq != do_deq;
  assign GEN_21 = T_1289 ? do_enq : maybe_full;
  assign T_1291 = T_1157 == 1'h0;
  assign T_1421 = 1'h0 - 1'h0;
  assign ptr_diff = T_1421[0:0];
  assign T_1423 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[1:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_4[2:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  GEN_6 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_a_type[initvar] = GEN_6[2:0];
  GEN_7 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_union[initvar] = GEN_7[11:0];
  GEN_8 = {2{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_8[63:0];
  GEN_9 = {1{$random}};
  maybe_full = GEN_9[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1160_en & ram_header_src_T_1160_mask) begin
      ram_header_src[ram_header_src_T_1160_addr] <= ram_header_src_T_1160_data;
    end
    if(ram_header_dst_T_1160_en & ram_header_dst_T_1160_mask) begin
      ram_header_dst[ram_header_dst_T_1160_addr] <= ram_header_dst_T_1160_data;
    end
    if(ram_payload_addr_block_T_1160_en & ram_payload_addr_block_T_1160_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1160_addr] <= ram_payload_addr_block_T_1160_data;
    end
    if(ram_payload_client_xact_id_T_1160_en & ram_payload_client_xact_id_T_1160_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1160_addr] <= ram_payload_client_xact_id_T_1160_data;
    end
    if(ram_payload_addr_beat_T_1160_en & ram_payload_addr_beat_T_1160_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1160_addr] <= ram_payload_addr_beat_T_1160_data;
    end
    if(ram_payload_is_builtin_type_T_1160_en & ram_payload_is_builtin_type_T_1160_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1160_addr] <= ram_payload_is_builtin_type_T_1160_data;
    end
    if(ram_payload_a_type_T_1160_en & ram_payload_a_type_T_1160_mask) begin
      ram_payload_a_type[ram_payload_a_type_T_1160_addr] <= ram_payload_a_type_T_1160_data;
    end
    if(ram_payload_union_T_1160_en & ram_payload_union_T_1160_mask) begin
      ram_payload_union[ram_payload_union_T_1160_addr] <= ram_payload_union_T_1160_data;
    end
    if(ram_payload_data_T_1160_en & ram_payload_data_T_1160_mask) begin
      ram_payload_data[ram_payload_data_T_1160_addr] <= ram_payload_data_T_1160_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1289) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_4(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_p_type,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_p_type,
  output  io_count
);
  reg [1:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1244_data;
  wire  ram_header_src_T_1244_addr;
  wire  ram_header_src_T_1244_en;
  wire [1:0] ram_header_src_T_1115_data;
  wire  ram_header_src_T_1115_addr;
  wire  ram_header_src_T_1115_mask;
  wire  ram_header_src_T_1115_en;
  reg [1:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1244_data;
  wire  ram_header_dst_T_1244_addr;
  wire  ram_header_dst_T_1244_en;
  wire [1:0] ram_header_dst_T_1115_data;
  wire  ram_header_dst_T_1115_addr;
  wire  ram_header_dst_T_1115_mask;
  wire  ram_header_dst_T_1115_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1244_data;
  wire  ram_payload_addr_block_T_1244_addr;
  wire  ram_payload_addr_block_T_1244_en;
  wire [25:0] ram_payload_addr_block_T_1115_data;
  wire  ram_payload_addr_block_T_1115_addr;
  wire  ram_payload_addr_block_T_1115_mask;
  wire  ram_payload_addr_block_T_1115_en;
  reg [1:0] ram_payload_p_type [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_p_type_T_1244_data;
  wire  ram_payload_p_type_T_1244_addr;
  wire  ram_payload_p_type_T_1244_en;
  wire [1:0] ram_payload_p_type_T_1115_data;
  wire  ram_payload_p_type_T_1115_addr;
  wire  ram_payload_p_type_T_1115_mask;
  wire  ram_payload_p_type_T_1115_en;
  reg  maybe_full;
  reg [31:0] GEN_4;
  wire  T_1112;
  wire  T_1113;
  wire  do_enq;
  wire  T_1114;
  wire  do_deq;
  wire  T_1239;
  wire  GEN_11;
  wire  T_1241;
  wire [1:0] T_1366;
  wire  ptr_diff;
  wire [1:0] T_1368;
  assign io_enq_ready = T_1112;
  assign io_deq_valid = T_1241;
  assign io_deq_bits_header_src = ram_header_src_T_1244_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1244_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1244_data;
  assign io_deq_bits_payload_p_type = ram_payload_p_type_T_1244_data;
  assign io_count = T_1368[0];
  assign ram_header_src_T_1244_addr = 1'h0;
  assign ram_header_src_T_1244_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_src_T_1244_data = ram_header_src[ram_header_src_T_1244_addr];
  `else
  assign ram_header_src_T_1244_data = ram_header_src_T_1244_addr >= 1'h1 ? $random : ram_header_src[ram_header_src_T_1244_addr];
  `endif
  assign ram_header_src_T_1115_data = io_enq_bits_header_src;
  assign ram_header_src_T_1115_addr = 1'h0;
  assign ram_header_src_T_1115_mask = do_enq;
  assign ram_header_src_T_1115_en = do_enq;
  assign ram_header_dst_T_1244_addr = 1'h0;
  assign ram_header_dst_T_1244_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_dst_T_1244_data = ram_header_dst[ram_header_dst_T_1244_addr];
  `else
  assign ram_header_dst_T_1244_data = ram_header_dst_T_1244_addr >= 1'h1 ? $random : ram_header_dst[ram_header_dst_T_1244_addr];
  `endif
  assign ram_header_dst_T_1115_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1115_addr = 1'h0;
  assign ram_header_dst_T_1115_mask = do_enq;
  assign ram_header_dst_T_1115_en = do_enq;
  assign ram_payload_addr_block_T_1244_addr = 1'h0;
  assign ram_payload_addr_block_T_1244_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_block_T_1244_data = ram_payload_addr_block[ram_payload_addr_block_T_1244_addr];
  `else
  assign ram_payload_addr_block_T_1244_data = ram_payload_addr_block_T_1244_addr >= 1'h1 ? $random : ram_payload_addr_block[ram_payload_addr_block_T_1244_addr];
  `endif
  assign ram_payload_addr_block_T_1115_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1115_addr = 1'h0;
  assign ram_payload_addr_block_T_1115_mask = do_enq;
  assign ram_payload_addr_block_T_1115_en = do_enq;
  assign ram_payload_p_type_T_1244_addr = 1'h0;
  assign ram_payload_p_type_T_1244_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_p_type_T_1244_data = ram_payload_p_type[ram_payload_p_type_T_1244_addr];
  `else
  assign ram_payload_p_type_T_1244_data = ram_payload_p_type_T_1244_addr >= 1'h1 ? $random : ram_payload_p_type[ram_payload_p_type_T_1244_addr];
  `endif
  assign ram_payload_p_type_T_1115_data = io_enq_bits_payload_p_type;
  assign ram_payload_p_type_T_1115_addr = 1'h0;
  assign ram_payload_p_type_T_1115_mask = do_enq;
  assign ram_payload_p_type_T_1115_en = do_enq;
  assign T_1112 = maybe_full == 1'h0;
  assign T_1113 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1113;
  assign T_1114 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1114;
  assign T_1239 = do_enq != do_deq;
  assign GEN_11 = T_1239 ? do_enq : maybe_full;
  assign T_1241 = T_1112 == 1'h0;
  assign T_1366 = 1'h0 - 1'h0;
  assign ptr_diff = T_1366[0:0];
  assign T_1368 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_p_type[initvar] = GEN_3[1:0];
  GEN_4 = {1{$random}};
  maybe_full = GEN_4[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1115_en & ram_header_src_T_1115_mask) begin
      ram_header_src[ram_header_src_T_1115_addr] <= ram_header_src_T_1115_data;
    end
    if(ram_header_dst_T_1115_en & ram_header_dst_T_1115_mask) begin
      ram_header_dst[ram_header_dst_T_1115_addr] <= ram_header_dst_T_1115_data;
    end
    if(ram_payload_addr_block_T_1115_en & ram_payload_addr_block_T_1115_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1115_addr] <= ram_payload_addr_block_T_1115_data;
    end
    if(ram_payload_p_type_T_1115_en & ram_payload_p_type_T_1115_mask) begin
      ram_payload_p_type[ram_payload_p_type_T_1115_addr] <= ram_payload_p_type_T_1115_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1239) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_5(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input   io_enq_bits_payload_voluntary,
  input  [2:0] io_enq_bits_payload_r_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output  io_deq_bits_payload_voluntary,
  output [2:0] io_deq_bits_payload_r_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [1:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1294_data;
  wire  ram_header_src_T_1294_addr;
  wire  ram_header_src_T_1294_en;
  wire [1:0] ram_header_src_T_1153_data;
  wire  ram_header_src_T_1153_addr;
  wire  ram_header_src_T_1153_mask;
  wire  ram_header_src_T_1153_en;
  reg [1:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1294_data;
  wire  ram_header_dst_T_1294_addr;
  wire  ram_header_dst_T_1294_en;
  wire [1:0] ram_header_dst_T_1153_data;
  wire  ram_header_dst_T_1153_addr;
  wire  ram_header_dst_T_1153_mask;
  wire  ram_header_dst_T_1153_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1294_data;
  wire  ram_payload_addr_beat_T_1294_addr;
  wire  ram_payload_addr_beat_T_1294_en;
  wire [2:0] ram_payload_addr_beat_T_1153_data;
  wire  ram_payload_addr_beat_T_1153_addr;
  wire  ram_payload_addr_beat_T_1153_mask;
  wire  ram_payload_addr_beat_T_1153_en;
  reg [25:0] ram_payload_addr_block [0:1];
  reg [31:0] GEN_3;
  wire [25:0] ram_payload_addr_block_T_1294_data;
  wire  ram_payload_addr_block_T_1294_addr;
  wire  ram_payload_addr_block_T_1294_en;
  wire [25:0] ram_payload_addr_block_T_1153_data;
  wire  ram_payload_addr_block_T_1153_addr;
  wire  ram_payload_addr_block_T_1153_mask;
  wire  ram_payload_addr_block_T_1153_en;
  reg [1:0] ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_4;
  wire [1:0] ram_payload_client_xact_id_T_1294_data;
  wire  ram_payload_client_xact_id_T_1294_addr;
  wire  ram_payload_client_xact_id_T_1294_en;
  wire [1:0] ram_payload_client_xact_id_T_1153_data;
  wire  ram_payload_client_xact_id_T_1153_addr;
  wire  ram_payload_client_xact_id_T_1153_mask;
  wire  ram_payload_client_xact_id_T_1153_en;
  reg  ram_payload_voluntary [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_voluntary_T_1294_data;
  wire  ram_payload_voluntary_T_1294_addr;
  wire  ram_payload_voluntary_T_1294_en;
  wire  ram_payload_voluntary_T_1153_data;
  wire  ram_payload_voluntary_T_1153_addr;
  wire  ram_payload_voluntary_T_1153_mask;
  wire  ram_payload_voluntary_T_1153_en;
  reg [2:0] ram_payload_r_type [0:1];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_r_type_T_1294_data;
  wire  ram_payload_r_type_T_1294_addr;
  wire  ram_payload_r_type_T_1294_en;
  wire [2:0] ram_payload_r_type_T_1153_data;
  wire  ram_payload_r_type_T_1153_addr;
  wire  ram_payload_r_type_T_1153_mask;
  wire  ram_payload_r_type_T_1153_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1294_data;
  wire  ram_payload_data_T_1294_addr;
  wire  ram_payload_data_T_1294_en;
  wire [63:0] ram_payload_data_T_1153_data;
  wire  ram_payload_data_T_1153_addr;
  wire  ram_payload_data_T_1153_mask;
  wire  ram_payload_data_T_1153_en;
  reg  T_1145;
  reg [31:0] GEN_8;
  reg  T_1147;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1150;
  wire  empty;
  wire  full;
  wire  T_1151;
  wire  do_enq;
  wire  T_1152;
  wire  do_deq;
  wire [1:0] T_1282;
  wire  T_1283;
  wire  GEN_19;
  wire [1:0] T_1287;
  wire  T_1288;
  wire  GEN_20;
  wire  T_1289;
  wire  GEN_21;
  wire  T_1291;
  wire  T_1293;
  wire [1:0] T_1420;
  wire  ptr_diff;
  wire  T_1421;
  wire [1:0] T_1422;
  assign io_enq_ready = T_1293;
  assign io_deq_valid = T_1291;
  assign io_deq_bits_header_src = ram_header_src_T_1294_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1294_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1294_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1294_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1294_data;
  assign io_deq_bits_payload_voluntary = ram_payload_voluntary_T_1294_data;
  assign io_deq_bits_payload_r_type = ram_payload_r_type_T_1294_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1294_data;
  assign io_count = T_1422;
  assign ram_header_src_T_1294_addr = T_1147;
  assign ram_header_src_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_src_T_1294_data = ram_header_src[ram_header_src_T_1294_addr];
  `else
  assign ram_header_src_T_1294_data = ram_header_src_T_1294_addr >= 2'h2 ? $random : ram_header_src[ram_header_src_T_1294_addr];
  `endif
  assign ram_header_src_T_1153_data = io_enq_bits_header_src;
  assign ram_header_src_T_1153_addr = T_1145;
  assign ram_header_src_T_1153_mask = do_enq;
  assign ram_header_src_T_1153_en = do_enq;
  assign ram_header_dst_T_1294_addr = T_1147;
  assign ram_header_dst_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_dst_T_1294_data = ram_header_dst[ram_header_dst_T_1294_addr];
  `else
  assign ram_header_dst_T_1294_data = ram_header_dst_T_1294_addr >= 2'h2 ? $random : ram_header_dst[ram_header_dst_T_1294_addr];
  `endif
  assign ram_header_dst_T_1153_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1153_addr = T_1145;
  assign ram_header_dst_T_1153_mask = do_enq;
  assign ram_header_dst_T_1153_en = do_enq;
  assign ram_payload_addr_beat_T_1294_addr = T_1147;
  assign ram_payload_addr_beat_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `else
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat_T_1294_addr >= 2'h2 ? $random : ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `endif
  assign ram_payload_addr_beat_T_1153_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1153_addr = T_1145;
  assign ram_payload_addr_beat_T_1153_mask = do_enq;
  assign ram_payload_addr_beat_T_1153_en = do_enq;
  assign ram_payload_addr_block_T_1294_addr = T_1147;
  assign ram_payload_addr_block_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_block_T_1294_data = ram_payload_addr_block[ram_payload_addr_block_T_1294_addr];
  `else
  assign ram_payload_addr_block_T_1294_data = ram_payload_addr_block_T_1294_addr >= 2'h2 ? $random : ram_payload_addr_block[ram_payload_addr_block_T_1294_addr];
  `endif
  assign ram_payload_addr_block_T_1153_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1153_addr = T_1145;
  assign ram_payload_addr_block_T_1153_mask = do_enq;
  assign ram_payload_addr_block_T_1153_en = do_enq;
  assign ram_payload_client_xact_id_T_1294_addr = T_1147;
  assign ram_payload_client_xact_id_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `else
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id_T_1294_addr >= 2'h2 ? $random : ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `endif
  assign ram_payload_client_xact_id_T_1153_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1153_addr = T_1145;
  assign ram_payload_client_xact_id_T_1153_mask = do_enq;
  assign ram_payload_client_xact_id_T_1153_en = do_enq;
  assign ram_payload_voluntary_T_1294_addr = T_1147;
  assign ram_payload_voluntary_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_voluntary_T_1294_data = ram_payload_voluntary[ram_payload_voluntary_T_1294_addr];
  `else
  assign ram_payload_voluntary_T_1294_data = ram_payload_voluntary_T_1294_addr >= 2'h2 ? $random : ram_payload_voluntary[ram_payload_voluntary_T_1294_addr];
  `endif
  assign ram_payload_voluntary_T_1153_data = io_enq_bits_payload_voluntary;
  assign ram_payload_voluntary_T_1153_addr = T_1145;
  assign ram_payload_voluntary_T_1153_mask = do_enq;
  assign ram_payload_voluntary_T_1153_en = do_enq;
  assign ram_payload_r_type_T_1294_addr = T_1147;
  assign ram_payload_r_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_r_type_T_1294_data = ram_payload_r_type[ram_payload_r_type_T_1294_addr];
  `else
  assign ram_payload_r_type_T_1294_data = ram_payload_r_type_T_1294_addr >= 2'h2 ? $random : ram_payload_r_type[ram_payload_r_type_T_1294_addr];
  `endif
  assign ram_payload_r_type_T_1153_data = io_enq_bits_payload_r_type;
  assign ram_payload_r_type_T_1153_addr = T_1145;
  assign ram_payload_r_type_T_1153_mask = do_enq;
  assign ram_payload_r_type_T_1153_en = do_enq;
  assign ram_payload_data_T_1294_addr = T_1147;
  assign ram_payload_data_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_data_T_1294_data = ram_payload_data[ram_payload_data_T_1294_addr];
  `else
  assign ram_payload_data_T_1294_data = ram_payload_data_T_1294_addr >= 2'h2 ? $random : ram_payload_data[ram_payload_data_T_1294_addr];
  `endif
  assign ram_payload_data_T_1153_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1153_addr = T_1145;
  assign ram_payload_data_T_1153_mask = do_enq;
  assign ram_payload_data_T_1153_en = do_enq;
  assign ptr_match = T_1145 == T_1147;
  assign T_1150 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1150;
  assign full = ptr_match & maybe_full;
  assign T_1151 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1151;
  assign T_1152 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1152;
  assign T_1282 = T_1145 + 1'h1;
  assign T_1283 = T_1282[0:0];
  assign GEN_19 = do_enq ? T_1283 : T_1145;
  assign T_1287 = T_1147 + 1'h1;
  assign T_1288 = T_1287[0:0];
  assign GEN_20 = do_deq ? T_1288 : T_1147;
  assign T_1289 = do_enq != do_deq;
  assign GEN_21 = T_1289 ? do_enq : maybe_full;
  assign T_1291 = empty == 1'h0;
  assign T_1293 = full == 1'h0;
  assign T_1420 = T_1145 - T_1147;
  assign ptr_diff = T_1420[0:0];
  assign T_1421 = maybe_full & ptr_match;
  assign T_1422 = {T_1421,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_3[25:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_4[1:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_voluntary[initvar] = GEN_5[0:0];
  GEN_6 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_r_type[initvar] = GEN_6[2:0];
  GEN_7 = {2{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  GEN_8 = {1{$random}};
  T_1145 = GEN_8[0:0];
  GEN_9 = {1{$random}};
  T_1147 = GEN_9[0:0];
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1153_en & ram_header_src_T_1153_mask) begin
      ram_header_src[ram_header_src_T_1153_addr] <= ram_header_src_T_1153_data;
    end
    if(ram_header_dst_T_1153_en & ram_header_dst_T_1153_mask) begin
      ram_header_dst[ram_header_dst_T_1153_addr] <= ram_header_dst_T_1153_data;
    end
    if(ram_payload_addr_beat_T_1153_en & ram_payload_addr_beat_T_1153_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1153_addr] <= ram_payload_addr_beat_T_1153_data;
    end
    if(ram_payload_addr_block_T_1153_en & ram_payload_addr_block_T_1153_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1153_addr] <= ram_payload_addr_block_T_1153_data;
    end
    if(ram_payload_client_xact_id_T_1153_en & ram_payload_client_xact_id_T_1153_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1153_addr] <= ram_payload_client_xact_id_T_1153_data;
    end
    if(ram_payload_voluntary_T_1153_en & ram_payload_voluntary_T_1153_mask) begin
      ram_payload_voluntary[ram_payload_voluntary_T_1153_addr] <= ram_payload_voluntary_T_1153_data;
    end
    if(ram_payload_r_type_T_1153_en & ram_payload_r_type_T_1153_mask) begin
      ram_payload_r_type[ram_payload_r_type_T_1153_addr] <= ram_payload_r_type_T_1153_data;
    end
    if(ram_payload_data_T_1153_en & ram_payload_data_T_1153_mask) begin
      ram_payload_data[ram_payload_data_T_1153_addr] <= ram_payload_data_T_1153_data;
    end
    if(reset) begin
      T_1145 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_1145 <= T_1283;
      end
    end
    if(reset) begin
      T_1147 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_1147 <= T_1288;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1289) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_6(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input  [2:0] io_enq_bits_payload_manager_xact_id,
  input   io_enq_bits_payload_is_builtin_type,
  input  [3:0] io_enq_bits_payload_g_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output [2:0] io_deq_bits_payload_manager_xact_id,
  output  io_deq_bits_payload_is_builtin_type,
  output [3:0] io_deq_bits_payload_g_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [1:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1294_data;
  wire  ram_header_src_T_1294_addr;
  wire  ram_header_src_T_1294_en;
  wire [1:0] ram_header_src_T_1153_data;
  wire  ram_header_src_T_1153_addr;
  wire  ram_header_src_T_1153_mask;
  wire  ram_header_src_T_1153_en;
  reg [1:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1294_data;
  wire  ram_header_dst_T_1294_addr;
  wire  ram_header_dst_T_1294_en;
  wire [1:0] ram_header_dst_T_1153_data;
  wire  ram_header_dst_T_1153_addr;
  wire  ram_header_dst_T_1153_mask;
  wire  ram_header_dst_T_1153_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1294_data;
  wire  ram_payload_addr_beat_T_1294_addr;
  wire  ram_payload_addr_beat_T_1294_en;
  wire [2:0] ram_payload_addr_beat_T_1153_data;
  wire  ram_payload_addr_beat_T_1153_addr;
  wire  ram_payload_addr_beat_T_1153_mask;
  wire  ram_payload_addr_beat_T_1153_en;
  reg [1:0] ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_client_xact_id_T_1294_data;
  wire  ram_payload_client_xact_id_T_1294_addr;
  wire  ram_payload_client_xact_id_T_1294_en;
  wire [1:0] ram_payload_client_xact_id_T_1153_data;
  wire  ram_payload_client_xact_id_T_1153_addr;
  wire  ram_payload_client_xact_id_T_1153_mask;
  wire  ram_payload_client_xact_id_T_1153_en;
  reg [2:0] ram_payload_manager_xact_id [0:1];
  reg [31:0] GEN_4;
  wire [2:0] ram_payload_manager_xact_id_T_1294_data;
  wire  ram_payload_manager_xact_id_T_1294_addr;
  wire  ram_payload_manager_xact_id_T_1294_en;
  wire [2:0] ram_payload_manager_xact_id_T_1153_data;
  wire  ram_payload_manager_xact_id_T_1153_addr;
  wire  ram_payload_manager_xact_id_T_1153_mask;
  wire  ram_payload_manager_xact_id_T_1153_en;
  reg  ram_payload_is_builtin_type [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1294_data;
  wire  ram_payload_is_builtin_type_T_1294_addr;
  wire  ram_payload_is_builtin_type_T_1294_en;
  wire  ram_payload_is_builtin_type_T_1153_data;
  wire  ram_payload_is_builtin_type_T_1153_addr;
  wire  ram_payload_is_builtin_type_T_1153_mask;
  wire  ram_payload_is_builtin_type_T_1153_en;
  reg [3:0] ram_payload_g_type [0:1];
  reg [31:0] GEN_6;
  wire [3:0] ram_payload_g_type_T_1294_data;
  wire  ram_payload_g_type_T_1294_addr;
  wire  ram_payload_g_type_T_1294_en;
  wire [3:0] ram_payload_g_type_T_1153_data;
  wire  ram_payload_g_type_T_1153_addr;
  wire  ram_payload_g_type_T_1153_mask;
  wire  ram_payload_g_type_T_1153_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1294_data;
  wire  ram_payload_data_T_1294_addr;
  wire  ram_payload_data_T_1294_en;
  wire [63:0] ram_payload_data_T_1153_data;
  wire  ram_payload_data_T_1153_addr;
  wire  ram_payload_data_T_1153_mask;
  wire  ram_payload_data_T_1153_en;
  reg  T_1145;
  reg [31:0] GEN_8;
  reg  T_1147;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1150;
  wire  empty;
  wire  full;
  wire  T_1151;
  wire  do_enq;
  wire  T_1152;
  wire  do_deq;
  wire [1:0] T_1282;
  wire  T_1283;
  wire  GEN_19;
  wire [1:0] T_1287;
  wire  T_1288;
  wire  GEN_20;
  wire  T_1289;
  wire  GEN_21;
  wire  T_1291;
  wire  T_1293;
  wire [1:0] T_1420;
  wire  ptr_diff;
  wire  T_1421;
  wire [1:0] T_1422;
  assign io_enq_ready = T_1293;
  assign io_deq_valid = T_1291;
  assign io_deq_bits_header_src = ram_header_src_T_1294_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1294_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1294_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1294_data;
  assign io_deq_bits_payload_manager_xact_id = ram_payload_manager_xact_id_T_1294_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1294_data;
  assign io_deq_bits_payload_g_type = ram_payload_g_type_T_1294_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1294_data;
  assign io_count = T_1422;
  assign ram_header_src_T_1294_addr = T_1147;
  assign ram_header_src_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_src_T_1294_data = ram_header_src[ram_header_src_T_1294_addr];
  `else
  assign ram_header_src_T_1294_data = ram_header_src_T_1294_addr >= 2'h2 ? $random : ram_header_src[ram_header_src_T_1294_addr];
  `endif
  assign ram_header_src_T_1153_data = io_enq_bits_header_src;
  assign ram_header_src_T_1153_addr = T_1145;
  assign ram_header_src_T_1153_mask = do_enq;
  assign ram_header_src_T_1153_en = do_enq;
  assign ram_header_dst_T_1294_addr = T_1147;
  assign ram_header_dst_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_dst_T_1294_data = ram_header_dst[ram_header_dst_T_1294_addr];
  `else
  assign ram_header_dst_T_1294_data = ram_header_dst_T_1294_addr >= 2'h2 ? $random : ram_header_dst[ram_header_dst_T_1294_addr];
  `endif
  assign ram_header_dst_T_1153_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1153_addr = T_1145;
  assign ram_header_dst_T_1153_mask = do_enq;
  assign ram_header_dst_T_1153_en = do_enq;
  assign ram_payload_addr_beat_T_1294_addr = T_1147;
  assign ram_payload_addr_beat_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `else
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat_T_1294_addr >= 2'h2 ? $random : ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `endif
  assign ram_payload_addr_beat_T_1153_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1153_addr = T_1145;
  assign ram_payload_addr_beat_T_1153_mask = do_enq;
  assign ram_payload_addr_beat_T_1153_en = do_enq;
  assign ram_payload_client_xact_id_T_1294_addr = T_1147;
  assign ram_payload_client_xact_id_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `else
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id_T_1294_addr >= 2'h2 ? $random : ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `endif
  assign ram_payload_client_xact_id_T_1153_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1153_addr = T_1145;
  assign ram_payload_client_xact_id_T_1153_mask = do_enq;
  assign ram_payload_client_xact_id_T_1153_en = do_enq;
  assign ram_payload_manager_xact_id_T_1294_addr = T_1147;
  assign ram_payload_manager_xact_id_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_manager_xact_id_T_1294_data = ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1294_addr];
  `else
  assign ram_payload_manager_xact_id_T_1294_data = ram_payload_manager_xact_id_T_1294_addr >= 2'h2 ? $random : ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1294_addr];
  `endif
  assign ram_payload_manager_xact_id_T_1153_data = io_enq_bits_payload_manager_xact_id;
  assign ram_payload_manager_xact_id_T_1153_addr = T_1145;
  assign ram_payload_manager_xact_id_T_1153_mask = do_enq;
  assign ram_payload_manager_xact_id_T_1153_en = do_enq;
  assign ram_payload_is_builtin_type_T_1294_addr = T_1147;
  assign ram_payload_is_builtin_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_is_builtin_type_T_1294_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1294_addr];
  `else
  assign ram_payload_is_builtin_type_T_1294_data = ram_payload_is_builtin_type_T_1294_addr >= 2'h2 ? $random : ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1294_addr];
  `endif
  assign ram_payload_is_builtin_type_T_1153_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1153_addr = T_1145;
  assign ram_payload_is_builtin_type_T_1153_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1153_en = do_enq;
  assign ram_payload_g_type_T_1294_addr = T_1147;
  assign ram_payload_g_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_g_type_T_1294_data = ram_payload_g_type[ram_payload_g_type_T_1294_addr];
  `else
  assign ram_payload_g_type_T_1294_data = ram_payload_g_type_T_1294_addr >= 2'h2 ? $random : ram_payload_g_type[ram_payload_g_type_T_1294_addr];
  `endif
  assign ram_payload_g_type_T_1153_data = io_enq_bits_payload_g_type;
  assign ram_payload_g_type_T_1153_addr = T_1145;
  assign ram_payload_g_type_T_1153_mask = do_enq;
  assign ram_payload_g_type_T_1153_en = do_enq;
  assign ram_payload_data_T_1294_addr = T_1147;
  assign ram_payload_data_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_data_T_1294_data = ram_payload_data[ram_payload_data_T_1294_addr];
  `else
  assign ram_payload_data_T_1294_data = ram_payload_data_T_1294_addr >= 2'h2 ? $random : ram_payload_data[ram_payload_data_T_1294_addr];
  `endif
  assign ram_payload_data_T_1153_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1153_addr = T_1145;
  assign ram_payload_data_T_1153_mask = do_enq;
  assign ram_payload_data_T_1153_en = do_enq;
  assign ptr_match = T_1145 == T_1147;
  assign T_1150 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1150;
  assign full = ptr_match & maybe_full;
  assign T_1151 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1151;
  assign T_1152 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1152;
  assign T_1282 = T_1145 + 1'h1;
  assign T_1283 = T_1282[0:0];
  assign GEN_19 = do_enq ? T_1283 : T_1145;
  assign T_1287 = T_1147 + 1'h1;
  assign T_1288 = T_1287[0:0];
  assign GEN_20 = do_deq ? T_1288 : T_1147;
  assign T_1289 = do_enq != do_deq;
  assign GEN_21 = T_1289 ? do_enq : maybe_full;
  assign T_1291 = empty == 1'h0;
  assign T_1293 = full == 1'h0;
  assign T_1420 = T_1145 - T_1147;
  assign ptr_diff = T_1420[0:0];
  assign T_1421 = maybe_full & ptr_match;
  assign T_1422 = {T_1421,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[1:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_manager_xact_id[initvar] = GEN_4[2:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  GEN_6 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_g_type[initvar] = GEN_6[3:0];
  GEN_7 = {2{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  GEN_8 = {1{$random}};
  T_1145 = GEN_8[0:0];
  GEN_9 = {1{$random}};
  T_1147 = GEN_9[0:0];
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1153_en & ram_header_src_T_1153_mask) begin
      ram_header_src[ram_header_src_T_1153_addr] <= ram_header_src_T_1153_data;
    end
    if(ram_header_dst_T_1153_en & ram_header_dst_T_1153_mask) begin
      ram_header_dst[ram_header_dst_T_1153_addr] <= ram_header_dst_T_1153_data;
    end
    if(ram_payload_addr_beat_T_1153_en & ram_payload_addr_beat_T_1153_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1153_addr] <= ram_payload_addr_beat_T_1153_data;
    end
    if(ram_payload_client_xact_id_T_1153_en & ram_payload_client_xact_id_T_1153_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1153_addr] <= ram_payload_client_xact_id_T_1153_data;
    end
    if(ram_payload_manager_xact_id_T_1153_en & ram_payload_manager_xact_id_T_1153_mask) begin
      ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1153_addr] <= ram_payload_manager_xact_id_T_1153_data;
    end
    if(ram_payload_is_builtin_type_T_1153_en & ram_payload_is_builtin_type_T_1153_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1153_addr] <= ram_payload_is_builtin_type_T_1153_data;
    end
    if(ram_payload_g_type_T_1153_en & ram_payload_g_type_T_1153_mask) begin
      ram_payload_g_type[ram_payload_g_type_T_1153_addr] <= ram_payload_g_type_T_1153_data;
    end
    if(ram_payload_data_T_1153_en & ram_payload_data_T_1153_mask) begin
      ram_payload_data[ram_payload_data_T_1153_addr] <= ram_payload_data_T_1153_data;
    end
    if(reset) begin
      T_1145 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_1145 <= T_1283;
      end
    end
    if(reset) begin
      T_1147 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_1147 <= T_1288;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1289) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module TileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_3_1_clk;
  wire  Queue_3_1_reset;
  wire  Queue_3_1_io_enq_ready;
  wire  Queue_3_1_io_enq_valid;
  wire [1:0] Queue_3_1_io_enq_bits_header_src;
  wire [1:0] Queue_3_1_io_enq_bits_header_dst;
  wire [25:0] Queue_3_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_3_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_3_1_io_enq_bits_payload_addr_beat;
  wire  Queue_3_1_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_3_1_io_enq_bits_payload_a_type;
  wire [11:0] Queue_3_1_io_enq_bits_payload_union;
  wire [63:0] Queue_3_1_io_enq_bits_payload_data;
  wire  Queue_3_1_io_deq_ready;
  wire  Queue_3_1_io_deq_valid;
  wire [1:0] Queue_3_1_io_deq_bits_header_src;
  wire [1:0] Queue_3_1_io_deq_bits_header_dst;
  wire [25:0] Queue_3_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_3_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_3_1_io_deq_bits_payload_addr_beat;
  wire  Queue_3_1_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_3_1_io_deq_bits_payload_a_type;
  wire [11:0] Queue_3_1_io_deq_bits_payload_union;
  wire [63:0] Queue_3_1_io_deq_bits_payload_data;
  wire  Queue_3_1_io_count;
  wire  Queue_4_1_clk;
  wire  Queue_4_1_reset;
  wire  Queue_4_1_io_enq_ready;
  wire  Queue_4_1_io_enq_valid;
  wire [1:0] Queue_4_1_io_enq_bits_header_src;
  wire [1:0] Queue_4_1_io_enq_bits_header_dst;
  wire [25:0] Queue_4_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_4_1_io_enq_bits_payload_p_type;
  wire  Queue_4_1_io_deq_ready;
  wire  Queue_4_1_io_deq_valid;
  wire [1:0] Queue_4_1_io_deq_bits_header_src;
  wire [1:0] Queue_4_1_io_deq_bits_header_dst;
  wire [25:0] Queue_4_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_4_1_io_deq_bits_payload_p_type;
  wire  Queue_4_1_io_count;
  wire  Queue_5_1_clk;
  wire  Queue_5_1_reset;
  wire  Queue_5_1_io_enq_ready;
  wire  Queue_5_1_io_enq_valid;
  wire [1:0] Queue_5_1_io_enq_bits_header_src;
  wire [1:0] Queue_5_1_io_enq_bits_header_dst;
  wire [2:0] Queue_5_1_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_5_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_5_1_io_enq_bits_payload_client_xact_id;
  wire  Queue_5_1_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_5_1_io_enq_bits_payload_r_type;
  wire [63:0] Queue_5_1_io_enq_bits_payload_data;
  wire  Queue_5_1_io_deq_ready;
  wire  Queue_5_1_io_deq_valid;
  wire [1:0] Queue_5_1_io_deq_bits_header_src;
  wire [1:0] Queue_5_1_io_deq_bits_header_dst;
  wire [2:0] Queue_5_1_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_5_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_5_1_io_deq_bits_payload_client_xact_id;
  wire  Queue_5_1_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_5_1_io_deq_bits_payload_r_type;
  wire [63:0] Queue_5_1_io_deq_bits_payload_data;
  wire [1:0] Queue_5_1_io_count;
  wire  Queue_6_1_clk;
  wire  Queue_6_1_reset;
  wire  Queue_6_1_io_enq_ready;
  wire  Queue_6_1_io_enq_valid;
  wire [1:0] Queue_6_1_io_enq_bits_header_src;
  wire [1:0] Queue_6_1_io_enq_bits_header_dst;
  wire [2:0] Queue_6_1_io_enq_bits_payload_addr_beat;
  wire [1:0] Queue_6_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_6_1_io_enq_bits_payload_manager_xact_id;
  wire  Queue_6_1_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_6_1_io_enq_bits_payload_g_type;
  wire [63:0] Queue_6_1_io_enq_bits_payload_data;
  wire  Queue_6_1_io_deq_ready;
  wire  Queue_6_1_io_deq_valid;
  wire [1:0] Queue_6_1_io_deq_bits_header_src;
  wire [1:0] Queue_6_1_io_deq_bits_header_dst;
  wire [2:0] Queue_6_1_io_deq_bits_payload_addr_beat;
  wire [1:0] Queue_6_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_6_1_io_deq_bits_payload_manager_xact_id;
  wire  Queue_6_1_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_6_1_io_deq_bits_payload_g_type;
  wire [63:0] Queue_6_1_io_deq_bits_payload_data;
  wire [1:0] Queue_6_1_io_count;
  Queue_3 Queue_3_1 (
    .clk(Queue_3_1_clk),
    .reset(Queue_3_1_reset),
    .io_enq_ready(Queue_3_1_io_enq_ready),
    .io_enq_valid(Queue_3_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_3_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_3_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_3_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_3_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_3_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_3_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_3_1_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_3_1_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_3_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_3_1_io_deq_ready),
    .io_deq_valid(Queue_3_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_3_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_3_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_3_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_3_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_3_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_3_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_3_1_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_3_1_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_3_1_io_deq_bits_payload_data),
    .io_count(Queue_3_1_io_count)
  );
  Queue_4 Queue_4_1 (
    .clk(Queue_4_1_clk),
    .reset(Queue_4_1_reset),
    .io_enq_ready(Queue_4_1_io_enq_ready),
    .io_enq_valid(Queue_4_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_4_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_4_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_4_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_4_1_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_4_1_io_deq_ready),
    .io_deq_valid(Queue_4_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_4_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_4_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_4_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_4_1_io_deq_bits_payload_p_type),
    .io_count(Queue_4_1_io_count)
  );
  Queue_5 Queue_5_1 (
    .clk(Queue_5_1_clk),
    .reset(Queue_5_1_reset),
    .io_enq_ready(Queue_5_1_io_enq_ready),
    .io_enq_valid(Queue_5_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_5_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_5_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_5_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_5_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_5_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_5_1_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_5_1_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_5_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_5_1_io_deq_ready),
    .io_deq_valid(Queue_5_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_5_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_5_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_5_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_5_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_5_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_5_1_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_5_1_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_5_1_io_deq_bits_payload_data),
    .io_count(Queue_5_1_io_count)
  );
  Queue_6 Queue_6_1 (
    .clk(Queue_6_1_clk),
    .reset(Queue_6_1_reset),
    .io_enq_ready(Queue_6_1_io_enq_ready),
    .io_enq_valid(Queue_6_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_6_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_6_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_6_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_6_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_6_1_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_6_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_6_1_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_6_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_6_1_io_deq_ready),
    .io_deq_valid(Queue_6_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_6_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_6_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_6_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_6_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_6_1_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_6_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_6_1_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_6_1_io_deq_bits_payload_data),
    .io_count(Queue_6_1_io_count)
  );
  assign io_client_acquire_ready = Queue_3_1_io_enq_ready;
  assign io_client_grant_valid = Queue_6_1_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_6_1_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_6_1_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_6_1_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_6_1_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_6_1_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_6_1_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_6_1_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_6_1_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_4_1_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_4_1_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_4_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_4_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_4_1_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_5_1_io_enq_ready;
  assign io_manager_acquire_valid = Queue_3_1_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_3_1_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_3_1_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_3_1_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_3_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_3_1_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_3_1_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_3_1_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_3_1_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_3_1_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_6_1_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_4_1_io_enq_ready;
  assign io_manager_release_valid = Queue_5_1_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_5_1_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_5_1_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_5_1_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_5_1_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_5_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_5_1_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_5_1_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_5_1_io_deq_bits_payload_data;
  assign Queue_3_1_clk = clk;
  assign Queue_3_1_reset = reset;
  assign Queue_3_1_io_enq_valid = io_client_acquire_valid;
  assign Queue_3_1_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_3_1_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_3_1_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_3_1_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_3_1_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_3_1_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_3_1_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_3_1_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_3_1_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_3_1_io_deq_ready = io_manager_acquire_ready;
  assign Queue_4_1_clk = clk;
  assign Queue_4_1_reset = reset;
  assign Queue_4_1_io_enq_valid = io_manager_probe_valid;
  assign Queue_4_1_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_4_1_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_4_1_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_4_1_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_4_1_io_deq_ready = io_client_probe_ready;
  assign Queue_5_1_clk = clk;
  assign Queue_5_1_reset = reset;
  assign Queue_5_1_io_enq_valid = io_client_release_valid;
  assign Queue_5_1_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_5_1_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_5_1_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_5_1_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_5_1_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_5_1_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_5_1_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_5_1_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_5_1_io_deq_ready = io_manager_release_ready;
  assign Queue_6_1_clk = clk;
  assign Queue_6_1_reset = reset;
  assign Queue_6_1_io_enq_valid = io_manager_grant_valid;
  assign Queue_6_1_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_6_1_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_6_1_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_6_1_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_6_1_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_6_1_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_6_1_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_6_1_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_6_1_io_deq_ready = io_client_grant_ready;
endmodule
module ClientTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input  [1:0] io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [11:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [25:0] io_client_probe_bits_addr_block,
  output [1:0] io_client_probe_bits_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_addr_beat,
  input  [25:0] io_client_release_bits_addr_block,
  input  [1:0] io_client_release_bits_client_xact_id,
  input   io_client_release_bits_voluntary,
  input  [2:0] io_client_release_bits_r_type,
  input  [63:0] io_client_release_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output [1:0] io_client_grant_bits_client_xact_id,
  output [2:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  output  io_client_grant_bits_manager_id,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [2:0] io_client_finish_bits_manager_xact_id,
  input   io_client_finish_bits_manager_id,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [1:0] io_network_acquire_bits_header_src,
  output [1:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output [1:0] io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [11:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [1:0] io_network_grant_bits_header_src,
  input  [1:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input  [1:0] io_network_grant_bits_payload_client_xact_id,
  input  [2:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [1:0] io_network_finish_bits_header_src,
  output [1:0] io_network_finish_bits_header_dst,
  output [2:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [1:0] io_network_probe_bits_header_src,
  input  [1:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [1:0] io_network_release_bits_header_src,
  output [1:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output [1:0] io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [1:0] acq_with_header_bits_header_src;
  wire [1:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire [1:0] acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [11:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_4395;
  wire  T_4397;
  wire  T_4403;
  wire  rel_with_header_ready;
  wire  rel_with_header_valid;
  wire [1:0] rel_with_header_bits_header_src;
  wire [1:0] rel_with_header_bits_header_dst;
  wire [2:0] rel_with_header_bits_payload_addr_beat;
  wire [25:0] rel_with_header_bits_payload_addr_block;
  wire [1:0] rel_with_header_bits_payload_client_xact_id;
  wire  rel_with_header_bits_payload_voluntary;
  wire [2:0] rel_with_header_bits_payload_r_type;
  wire [63:0] rel_with_header_bits_payload_data;
  wire [31:0] GEN_1;
  wire [31:0] T_5040;
  wire  T_5042;
  wire  T_5048;
  wire  fin_with_header_ready;
  wire  fin_with_header_valid;
  wire [1:0] fin_with_header_bits_header_src;
  wire [1:0] fin_with_header_bits_header_dst;
  wire [2:0] fin_with_header_bits_payload_manager_xact_id;
  wire  fin_with_header_bits_payload_manager_id;
  wire  prb_without_header_ready;
  wire  prb_without_header_valid;
  wire [25:0] prb_without_header_bits_addr_block;
  wire [1:0] prb_without_header_bits_p_type;
  wire  gnt_without_header_ready;
  wire  gnt_without_header_valid;
  wire [2:0] gnt_without_header_bits_addr_beat;
  wire [1:0] gnt_without_header_bits_client_xact_id;
  wire [2:0] gnt_without_header_bits_manager_xact_id;
  wire  gnt_without_header_bits_is_builtin_type;
  wire [3:0] gnt_without_header_bits_g_type;
  wire [63:0] gnt_without_header_bits_data;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_probe_valid = prb_without_header_valid;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign io_client_release_ready = rel_with_header_ready;
  assign io_client_grant_valid = gnt_without_header_valid;
  assign io_client_grant_bits_addr_beat = gnt_without_header_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = gnt_without_header_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = gnt_without_header_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = gnt_without_header_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = gnt_without_header_bits_g_type;
  assign io_client_grant_bits_data = gnt_without_header_bits_data;
  assign io_client_grant_bits_manager_id = io_network_grant_bits_header_src[0];
  assign io_client_finish_ready = fin_with_header_ready;
  assign io_network_acquire_valid = acq_with_header_valid;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = gnt_without_header_ready;
  assign io_network_finish_valid = fin_with_header_valid;
  assign io_network_finish_bits_header_src = fin_with_header_bits_header_src;
  assign io_network_finish_bits_header_dst = fin_with_header_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = fin_with_header_bits_payload_manager_xact_id;
  assign io_network_probe_ready = prb_without_header_ready;
  assign io_network_release_valid = rel_with_header_valid;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign acq_with_header_ready = io_network_acquire_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = {{1'd0}, 1'h0};
  assign acq_with_header_bits_header_dst = {{1'd0}, T_4403};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_4395 = GEN_0 << 6;
  assign T_4397 = 32'h80000000 <= T_4395;
  assign T_4403 = T_4397 ? 1'h0 : 1'h1;
  assign rel_with_header_ready = io_network_release_ready;
  assign rel_with_header_valid = io_client_release_valid;
  assign rel_with_header_bits_header_src = {{1'd0}, 1'h0};
  assign rel_with_header_bits_header_dst = {{1'd0}, T_5048};
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign GEN_1 = {{6'd0}, io_client_release_bits_addr_block};
  assign T_5040 = GEN_1 << 6;
  assign T_5042 = 32'h80000000 <= T_5040;
  assign T_5048 = T_5042 ? 1'h0 : 1'h1;
  assign fin_with_header_ready = io_network_finish_ready;
  assign fin_with_header_valid = io_client_finish_valid;
  assign fin_with_header_bits_header_src = {{1'd0}, 1'h0};
  assign fin_with_header_bits_header_dst = {{1'd0}, io_client_finish_bits_manager_id};
  assign fin_with_header_bits_payload_manager_xact_id = io_client_finish_bits_manager_xact_id;
  assign fin_with_header_bits_payload_manager_id = io_client_finish_bits_manager_id;
  assign prb_without_header_ready = io_client_probe_ready;
  assign prb_without_header_valid = io_network_probe_valid;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign gnt_without_header_ready = io_client_grant_ready;
  assign gnt_without_header_valid = io_network_grant_valid;
  assign gnt_without_header_bits_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign gnt_without_header_bits_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign gnt_without_header_bits_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign gnt_without_header_bits_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign gnt_without_header_bits_g_type = io_network_grant_bits_payload_g_type;
  assign gnt_without_header_bits_data = io_network_grant_bits_payload_data;
endmodule
module TileLinkEnqueuer_1(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_7_1_clk;
  wire  Queue_7_1_reset;
  wire  Queue_7_1_io_enq_ready;
  wire  Queue_7_1_io_enq_valid;
  wire [1:0] Queue_7_1_io_enq_bits_header_src;
  wire [1:0] Queue_7_1_io_enq_bits_header_dst;
  wire [25:0] Queue_7_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_7_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_7_1_io_enq_bits_payload_addr_beat;
  wire  Queue_7_1_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_7_1_io_enq_bits_payload_a_type;
  wire [11:0] Queue_7_1_io_enq_bits_payload_union;
  wire [63:0] Queue_7_1_io_enq_bits_payload_data;
  wire  Queue_7_1_io_deq_ready;
  wire  Queue_7_1_io_deq_valid;
  wire [1:0] Queue_7_1_io_deq_bits_header_src;
  wire [1:0] Queue_7_1_io_deq_bits_header_dst;
  wire [25:0] Queue_7_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_7_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_7_1_io_deq_bits_payload_addr_beat;
  wire  Queue_7_1_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_7_1_io_deq_bits_payload_a_type;
  wire [11:0] Queue_7_1_io_deq_bits_payload_union;
  wire [63:0] Queue_7_1_io_deq_bits_payload_data;
  wire  Queue_7_1_io_count;
  wire  Queue_8_1_clk;
  wire  Queue_8_1_reset;
  wire  Queue_8_1_io_enq_ready;
  wire  Queue_8_1_io_enq_valid;
  wire [1:0] Queue_8_1_io_enq_bits_header_src;
  wire [1:0] Queue_8_1_io_enq_bits_header_dst;
  wire [25:0] Queue_8_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_8_1_io_enq_bits_payload_p_type;
  wire  Queue_8_1_io_deq_ready;
  wire  Queue_8_1_io_deq_valid;
  wire [1:0] Queue_8_1_io_deq_bits_header_src;
  wire [1:0] Queue_8_1_io_deq_bits_header_dst;
  wire [25:0] Queue_8_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_8_1_io_deq_bits_payload_p_type;
  wire  Queue_8_1_io_count;
  wire  Queue_9_1_clk;
  wire  Queue_9_1_reset;
  wire  Queue_9_1_io_enq_ready;
  wire  Queue_9_1_io_enq_valid;
  wire [1:0] Queue_9_1_io_enq_bits_header_src;
  wire [1:0] Queue_9_1_io_enq_bits_header_dst;
  wire [2:0] Queue_9_1_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_9_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_9_1_io_enq_bits_payload_client_xact_id;
  wire  Queue_9_1_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_9_1_io_enq_bits_payload_r_type;
  wire [63:0] Queue_9_1_io_enq_bits_payload_data;
  wire  Queue_9_1_io_deq_ready;
  wire  Queue_9_1_io_deq_valid;
  wire [1:0] Queue_9_1_io_deq_bits_header_src;
  wire [1:0] Queue_9_1_io_deq_bits_header_dst;
  wire [2:0] Queue_9_1_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_9_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_9_1_io_deq_bits_payload_client_xact_id;
  wire  Queue_9_1_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_9_1_io_deq_bits_payload_r_type;
  wire [63:0] Queue_9_1_io_deq_bits_payload_data;
  wire [1:0] Queue_9_1_io_count;
  wire  Queue_10_1_clk;
  wire  Queue_10_1_reset;
  wire  Queue_10_1_io_enq_ready;
  wire  Queue_10_1_io_enq_valid;
  wire [1:0] Queue_10_1_io_enq_bits_header_src;
  wire [1:0] Queue_10_1_io_enq_bits_header_dst;
  wire [2:0] Queue_10_1_io_enq_bits_payload_addr_beat;
  wire [1:0] Queue_10_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_10_1_io_enq_bits_payload_manager_xact_id;
  wire  Queue_10_1_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_10_1_io_enq_bits_payload_g_type;
  wire [63:0] Queue_10_1_io_enq_bits_payload_data;
  wire  Queue_10_1_io_deq_ready;
  wire  Queue_10_1_io_deq_valid;
  wire [1:0] Queue_10_1_io_deq_bits_header_src;
  wire [1:0] Queue_10_1_io_deq_bits_header_dst;
  wire [2:0] Queue_10_1_io_deq_bits_payload_addr_beat;
  wire [1:0] Queue_10_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_10_1_io_deq_bits_payload_manager_xact_id;
  wire  Queue_10_1_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_10_1_io_deq_bits_payload_g_type;
  wire [63:0] Queue_10_1_io_deq_bits_payload_data;
  wire [1:0] Queue_10_1_io_count;
  Queue_3 Queue_7_1 (
    .clk(Queue_7_1_clk),
    .reset(Queue_7_1_reset),
    .io_enq_ready(Queue_7_1_io_enq_ready),
    .io_enq_valid(Queue_7_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_7_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_7_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_7_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_7_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_7_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_7_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_7_1_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_7_1_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_7_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_7_1_io_deq_ready),
    .io_deq_valid(Queue_7_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_7_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_7_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_7_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_7_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_7_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_7_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_7_1_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_7_1_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_7_1_io_deq_bits_payload_data),
    .io_count(Queue_7_1_io_count)
  );
  Queue_4 Queue_8_1 (
    .clk(Queue_8_1_clk),
    .reset(Queue_8_1_reset),
    .io_enq_ready(Queue_8_1_io_enq_ready),
    .io_enq_valid(Queue_8_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_8_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_8_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_8_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_8_1_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_8_1_io_deq_ready),
    .io_deq_valid(Queue_8_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_8_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_8_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_8_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_8_1_io_deq_bits_payload_p_type),
    .io_count(Queue_8_1_io_count)
  );
  Queue_5 Queue_9_1 (
    .clk(Queue_9_1_clk),
    .reset(Queue_9_1_reset),
    .io_enq_ready(Queue_9_1_io_enq_ready),
    .io_enq_valid(Queue_9_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_9_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_9_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_9_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_9_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_9_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_9_1_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_9_1_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_9_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_9_1_io_deq_ready),
    .io_deq_valid(Queue_9_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_9_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_9_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_9_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_9_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_9_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_9_1_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_9_1_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_9_1_io_deq_bits_payload_data),
    .io_count(Queue_9_1_io_count)
  );
  Queue_6 Queue_10_1 (
    .clk(Queue_10_1_clk),
    .reset(Queue_10_1_reset),
    .io_enq_ready(Queue_10_1_io_enq_ready),
    .io_enq_valid(Queue_10_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_10_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_10_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_10_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_10_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_10_1_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_10_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_10_1_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_10_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_10_1_io_deq_ready),
    .io_deq_valid(Queue_10_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_10_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_10_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_10_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_10_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_10_1_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_10_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_10_1_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_10_1_io_deq_bits_payload_data),
    .io_count(Queue_10_1_io_count)
  );
  assign io_client_acquire_ready = Queue_7_1_io_enq_ready;
  assign io_client_grant_valid = Queue_10_1_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_10_1_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_10_1_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_10_1_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_10_1_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_10_1_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_10_1_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_10_1_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_10_1_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_8_1_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_8_1_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_8_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_8_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_8_1_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_9_1_io_enq_ready;
  assign io_manager_acquire_valid = Queue_7_1_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_7_1_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_7_1_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_7_1_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_7_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_7_1_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_7_1_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_7_1_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_7_1_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_7_1_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_10_1_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_8_1_io_enq_ready;
  assign io_manager_release_valid = Queue_9_1_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_9_1_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_9_1_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_9_1_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_9_1_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_9_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_9_1_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_9_1_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_9_1_io_deq_bits_payload_data;
  assign Queue_7_1_clk = clk;
  assign Queue_7_1_reset = reset;
  assign Queue_7_1_io_enq_valid = io_client_acquire_valid;
  assign Queue_7_1_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_7_1_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_7_1_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_7_1_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_7_1_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_7_1_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_7_1_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_7_1_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_7_1_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_7_1_io_deq_ready = io_manager_acquire_ready;
  assign Queue_8_1_clk = clk;
  assign Queue_8_1_reset = reset;
  assign Queue_8_1_io_enq_valid = io_manager_probe_valid;
  assign Queue_8_1_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_8_1_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_8_1_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_8_1_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_8_1_io_deq_ready = io_client_probe_ready;
  assign Queue_9_1_clk = clk;
  assign Queue_9_1_reset = reset;
  assign Queue_9_1_io_enq_valid = io_client_release_valid;
  assign Queue_9_1_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_9_1_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_9_1_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_9_1_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_9_1_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_9_1_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_9_1_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_9_1_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_9_1_io_deq_ready = io_manager_release_ready;
  assign Queue_10_1_clk = clk;
  assign Queue_10_1_reset = reset;
  assign Queue_10_1_io_enq_valid = io_manager_grant_valid;
  assign Queue_10_1_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_10_1_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_10_1_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_10_1_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_10_1_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_10_1_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_10_1_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_10_1_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_10_1_io_deq_ready = io_client_grant_ready;
endmodule
module FinishQueue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output [1:0] io_count
);
  reg [2:0] T_244_manager_xact_id [0:1];
  reg [31:0] GEN_0;
  wire [2:0] T_244_manager_xact_id_T_301_data;
  wire  T_244_manager_xact_id_T_301_addr;
  wire  T_244_manager_xact_id_T_301_en;
  wire [2:0] T_244_manager_xact_id_T_260_data;
  wire  T_244_manager_xact_id_T_260_addr;
  wire  T_244_manager_xact_id_T_260_mask;
  wire  T_244_manager_xact_id_T_260_en;
  reg  T_244_manager_id [0:1];
  reg [31:0] GEN_1;
  wire  T_244_manager_id_T_301_data;
  wire  T_244_manager_id_T_301_addr;
  wire  T_244_manager_id_T_301_en;
  wire  T_244_manager_id_T_260_data;
  wire  T_244_manager_id_T_260_addr;
  wire  T_244_manager_id_T_260_mask;
  wire  T_244_manager_id_T_260_en;
  reg  T_246;
  reg [31:0] GEN_2;
  reg  T_248;
  reg [31:0] GEN_3;
  reg  T_250;
  reg [31:0] GEN_4;
  wire  T_251;
  wire  T_253;
  wire  T_254;
  wire  T_255;
  wire  T_256;
  wire  T_257;
  wire  T_258;
  wire  T_259;
  wire [1:0] T_289;
  wire  T_290;
  wire  GEN_7;
  wire [1:0] T_294;
  wire  T_295;
  wire  GEN_8;
  wire  T_296;
  wire  GEN_9;
  wire  T_298;
  wire  T_300;
  wire [1:0] T_327;
  wire  T_328;
  wire  T_329;
  wire [1:0] T_330;
  assign io_enq_ready = T_300;
  assign io_deq_valid = T_298;
  assign io_deq_bits_manager_xact_id = T_244_manager_xact_id_T_301_data;
  assign io_deq_bits_manager_id = T_244_manager_id_T_301_data;
  assign io_count = T_330;
  assign T_244_manager_xact_id_T_301_addr = T_248;
  assign T_244_manager_xact_id_T_301_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_244_manager_xact_id_T_301_data = T_244_manager_xact_id[T_244_manager_xact_id_T_301_addr];
  `else
  assign T_244_manager_xact_id_T_301_data = T_244_manager_xact_id_T_301_addr >= 2'h2 ? $random : T_244_manager_xact_id[T_244_manager_xact_id_T_301_addr];
  `endif
  assign T_244_manager_xact_id_T_260_data = io_enq_bits_manager_xact_id;
  assign T_244_manager_xact_id_T_260_addr = T_246;
  assign T_244_manager_xact_id_T_260_mask = T_257;
  assign T_244_manager_xact_id_T_260_en = T_257;
  assign T_244_manager_id_T_301_addr = T_248;
  assign T_244_manager_id_T_301_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_244_manager_id_T_301_data = T_244_manager_id[T_244_manager_id_T_301_addr];
  `else
  assign T_244_manager_id_T_301_data = T_244_manager_id_T_301_addr >= 2'h2 ? $random : T_244_manager_id[T_244_manager_id_T_301_addr];
  `endif
  assign T_244_manager_id_T_260_data = io_enq_bits_manager_id;
  assign T_244_manager_id_T_260_addr = T_246;
  assign T_244_manager_id_T_260_mask = T_257;
  assign T_244_manager_id_T_260_en = T_257;
  assign T_251 = T_246 == T_248;
  assign T_253 = T_250 == 1'h0;
  assign T_254 = T_251 & T_253;
  assign T_255 = T_251 & T_250;
  assign T_256 = io_enq_ready & io_enq_valid;
  assign T_257 = T_256;
  assign T_258 = io_deq_ready & io_deq_valid;
  assign T_259 = T_258;
  assign T_289 = T_246 + 1'h1;
  assign T_290 = T_289[0:0];
  assign GEN_7 = T_257 ? T_290 : T_246;
  assign T_294 = T_248 + 1'h1;
  assign T_295 = T_294[0:0];
  assign GEN_8 = T_259 ? T_295 : T_248;
  assign T_296 = T_257 != T_259;
  assign GEN_9 = T_296 ? T_257 : T_250;
  assign T_298 = T_254 == 1'h0;
  assign T_300 = T_255 == 1'h0;
  assign T_327 = T_246 - T_248;
  assign T_328 = T_327[0:0];
  assign T_329 = T_250 & T_251;
  assign T_330 = {T_329,T_328};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    T_244_manager_xact_id[initvar] = GEN_0[2:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    T_244_manager_id[initvar] = GEN_1[0:0];
  GEN_2 = {1{$random}};
  T_246 = GEN_2[0:0];
  GEN_3 = {1{$random}};
  T_248 = GEN_3[0:0];
  GEN_4 = {1{$random}};
  T_250 = GEN_4[0:0];
  end
`endif
  always @(posedge clk) begin
    if(T_244_manager_xact_id_T_260_en & T_244_manager_xact_id_T_260_mask) begin
      T_244_manager_xact_id[T_244_manager_xact_id_T_260_addr] <= T_244_manager_xact_id_T_260_data;
    end
    if(T_244_manager_id_T_260_en & T_244_manager_id_T_260_mask) begin
      T_244_manager_id[T_244_manager_id_T_260_addr] <= T_244_manager_id_T_260_data;
    end
    if(reset) begin
      T_246 <= 1'h0;
    end else begin
      if(T_257) begin
        T_246 <= T_290;
      end
    end
    if(reset) begin
      T_248 <= 1'h0;
    end else begin
      if(T_259) begin
        T_248 <= T_295;
      end
    end
    if(reset) begin
      T_250 <= 1'h0;
    end else begin
      if(T_296) begin
        T_250 <= T_257;
      end
    end
  end
endmodule
module FinishUnit(
  input   clk,
  input   reset,
  output  io_grant_ready,
  input   io_grant_valid,
  input  [1:0] io_grant_bits_header_src,
  input  [1:0] io_grant_bits_header_dst,
  input  [2:0] io_grant_bits_payload_addr_beat,
  input  [1:0] io_grant_bits_payload_client_xact_id,
  input  [2:0] io_grant_bits_payload_manager_xact_id,
  input   io_grant_bits_payload_is_builtin_type,
  input  [3:0] io_grant_bits_payload_g_type,
  input  [63:0] io_grant_bits_payload_data,
  input   io_refill_ready,
  output  io_refill_valid,
  output [2:0] io_refill_bits_addr_beat,
  output [1:0] io_refill_bits_client_xact_id,
  output [2:0] io_refill_bits_manager_xact_id,
  output  io_refill_bits_is_builtin_type,
  output [3:0] io_refill_bits_g_type,
  output [63:0] io_refill_bits_data,
  input   io_finish_ready,
  output  io_finish_valid,
  output [1:0] io_finish_bits_header_src,
  output [1:0] io_finish_bits_header_dst,
  output [2:0] io_finish_bits_payload_manager_xact_id,
  output  io_ready
);
  wire  T_1173;
  wire [2:0] T_1182_0;
  wire [3:0] GEN_1;
  wire  T_1184;
  wire [1:0] T_1192_0;
  wire [1:0] T_1192_1;
  wire [3:0] GEN_2;
  wire  T_1194;
  wire [3:0] GEN_3;
  wire  T_1195;
  wire  T_1198;
  wire  T_1199;
  wire  T_1201;
  reg [2:0] T_1203;
  reg [31:0] GEN_9;
  wire  T_1205;
  wire [2:0] GEN_4;
  wire [3:0] T_1207;
  wire [2:0] T_1208;
  wire [2:0] GEN_0;
  wire  T_1209;
  wire  T_1211;
  wire  FinishQueue_3_1_clk;
  wire  FinishQueue_3_1_reset;
  wire  FinishQueue_3_1_io_enq_ready;
  wire  FinishQueue_3_1_io_enq_valid;
  wire [2:0] FinishQueue_3_1_io_enq_bits_manager_xact_id;
  wire  FinishQueue_3_1_io_enq_bits_manager_id;
  wire  FinishQueue_3_1_io_deq_ready;
  wire  FinishQueue_3_1_io_deq_valid;
  wire [2:0] FinishQueue_3_1_io_deq_bits_manager_xact_id;
  wire  FinishQueue_3_1_io_deq_bits_manager_id;
  wire [1:0] FinishQueue_3_1_io_count;
  wire [3:0] GEN_5;
  wire  T_1243;
  wire  T_1244;
  wire  T_1246;
  wire  T_1248;
  wire [2:0] T_1256_0;
  wire [3:0] GEN_6;
  wire  T_1258;
  wire [1:0] T_1266_0;
  wire [1:0] T_1266_1;
  wire [3:0] GEN_7;
  wire  T_1268;
  wire [3:0] GEN_8;
  wire  T_1269;
  wire  T_1272;
  wire  T_1273;
  wire  T_1276;
  wire  T_1277;
  wire  T_1278;
  wire [2:0] T_1304_manager_xact_id;
  wire  T_1340;
  wire  T_1341;
  wire  T_1342;
  wire  T_1355;
  FinishQueue_3 FinishQueue_3_1 (
    .clk(FinishQueue_3_1_clk),
    .reset(FinishQueue_3_1_reset),
    .io_enq_ready(FinishQueue_3_1_io_enq_ready),
    .io_enq_valid(FinishQueue_3_1_io_enq_valid),
    .io_enq_bits_manager_xact_id(FinishQueue_3_1_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(FinishQueue_3_1_io_enq_bits_manager_id),
    .io_deq_ready(FinishQueue_3_1_io_deq_ready),
    .io_deq_valid(FinishQueue_3_1_io_deq_valid),
    .io_deq_bits_manager_xact_id(FinishQueue_3_1_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(FinishQueue_3_1_io_deq_bits_manager_id),
    .io_count(FinishQueue_3_1_io_count)
  );
  assign io_grant_ready = T_1355;
  assign io_refill_valid = T_1342;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_finish_valid = FinishQueue_3_1_io_deq_valid;
  assign io_finish_bits_header_src = {{1'd0}, 1'h1};
  assign io_finish_bits_header_dst = {{1'd0}, FinishQueue_3_1_io_deq_bits_manager_id};
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_3_1_io_deq_bits_manager_xact_id;
  assign io_ready = FinishQueue_3_1_io_enq_ready;
  assign T_1173 = io_grant_ready & io_grant_valid;
  assign T_1182_0 = 3'h5;
  assign GEN_1 = {{1'd0}, T_1182_0};
  assign T_1184 = GEN_1 == io_grant_bits_payload_g_type;
  assign T_1192_0 = 2'h0;
  assign T_1192_1 = 2'h1;
  assign GEN_2 = {{2'd0}, T_1192_0};
  assign T_1194 = GEN_2 == io_grant_bits_payload_g_type;
  assign GEN_3 = {{2'd0}, T_1192_1};
  assign T_1195 = GEN_3 == io_grant_bits_payload_g_type;
  assign T_1198 = T_1194 | T_1195;
  assign T_1199 = io_grant_bits_payload_is_builtin_type ? T_1184 : T_1198;
  assign T_1201 = T_1173 & T_1199;
  assign T_1205 = T_1203 == 3'h7;
  assign GEN_4 = {{2'd0}, 1'h1};
  assign T_1207 = T_1203 + GEN_4;
  assign T_1208 = T_1207[2:0];
  assign GEN_0 = T_1201 ? T_1208 : T_1203;
  assign T_1209 = T_1201 & T_1205;
  assign T_1211 = T_1199 ? T_1209 : T_1173;
  assign FinishQueue_3_1_clk = clk;
  assign FinishQueue_3_1_reset = reset;
  assign FinishQueue_3_1_io_enq_valid = T_1278;
  assign FinishQueue_3_1_io_enq_bits_manager_xact_id = T_1304_manager_xact_id;
  assign FinishQueue_3_1_io_enq_bits_manager_id = io_grant_bits_header_src[0];
  assign FinishQueue_3_1_io_deq_ready = io_finish_ready;
  assign GEN_5 = {{1'd0}, 3'h0};
  assign T_1243 = io_grant_bits_payload_g_type == GEN_5;
  assign T_1244 = io_grant_bits_payload_is_builtin_type & T_1243;
  assign T_1246 = T_1244 == 1'h0;
  assign T_1248 = T_1173 & T_1246;
  assign T_1256_0 = 3'h5;
  assign GEN_6 = {{1'd0}, T_1256_0};
  assign T_1258 = GEN_6 == io_grant_bits_payload_g_type;
  assign T_1266_0 = 2'h0;
  assign T_1266_1 = 2'h1;
  assign GEN_7 = {{2'd0}, T_1266_0};
  assign T_1268 = GEN_7 == io_grant_bits_payload_g_type;
  assign GEN_8 = {{2'd0}, T_1266_1};
  assign T_1269 = GEN_8 == io_grant_bits_payload_g_type;
  assign T_1272 = T_1268 | T_1269;
  assign T_1273 = io_grant_bits_payload_is_builtin_type ? T_1258 : T_1272;
  assign T_1276 = T_1273 == 1'h0;
  assign T_1277 = T_1276 | T_1211;
  assign T_1278 = T_1248 & T_1277;
  assign T_1304_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign T_1340 = T_1246 == 1'h0;
  assign T_1341 = FinishQueue_3_1_io_enq_ready | T_1340;
  assign T_1342 = T_1341 & io_grant_valid;
  assign T_1355 = T_1341 & io_refill_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  T_1203 = GEN_9[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1203 <= 3'h0;
    end else begin
      if(T_1201) begin
        T_1203 <= T_1208;
      end
    end
  end
endmodule
module ClientUncachedTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input  [1:0] io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [11:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output [1:0] io_client_grant_bits_client_xact_id,
  output [2:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [1:0] io_network_acquire_bits_header_src,
  output [1:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output [1:0] io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [11:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [1:0] io_network_grant_bits_header_src,
  input  [1:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input  [1:0] io_network_grant_bits_payload_client_xact_id,
  input  [2:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [1:0] io_network_finish_bits_header_src,
  output [1:0] io_network_finish_bits_header_dst,
  output [2:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [1:0] io_network_probe_bits_header_src,
  input  [1:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [1:0] io_network_release_bits_header_src,
  output [1:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output [1:0] io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  finisher_clk;
  wire  finisher_reset;
  wire  finisher_io_grant_ready;
  wire  finisher_io_grant_valid;
  wire [1:0] finisher_io_grant_bits_header_src;
  wire [1:0] finisher_io_grant_bits_header_dst;
  wire [2:0] finisher_io_grant_bits_payload_addr_beat;
  wire [1:0] finisher_io_grant_bits_payload_client_xact_id;
  wire [2:0] finisher_io_grant_bits_payload_manager_xact_id;
  wire  finisher_io_grant_bits_payload_is_builtin_type;
  wire [3:0] finisher_io_grant_bits_payload_g_type;
  wire [63:0] finisher_io_grant_bits_payload_data;
  wire  finisher_io_refill_ready;
  wire  finisher_io_refill_valid;
  wire [2:0] finisher_io_refill_bits_addr_beat;
  wire [1:0] finisher_io_refill_bits_client_xact_id;
  wire [2:0] finisher_io_refill_bits_manager_xact_id;
  wire  finisher_io_refill_bits_is_builtin_type;
  wire [3:0] finisher_io_refill_bits_g_type;
  wire [63:0] finisher_io_refill_bits_data;
  wire  finisher_io_finish_ready;
  wire  finisher_io_finish_valid;
  wire [1:0] finisher_io_finish_bits_header_src;
  wire [1:0] finisher_io_finish_bits_header_dst;
  wire [2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire  finisher_io_ready;
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [1:0] acq_with_header_bits_header_src;
  wire [1:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire [1:0] acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [11:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3765;
  wire  T_3767;
  wire  T_3773;
  wire  T_3774;
  wire  T_3775;
  reg [1:0] GEN_1;
  reg [31:0] GEN_9;
  reg [1:0] GEN_2;
  reg [31:0] GEN_10;
  reg [2:0] GEN_3;
  reg [31:0] GEN_11;
  reg [25:0] GEN_4;
  reg [31:0] GEN_12;
  reg [1:0] GEN_5;
  reg [31:0] GEN_13;
  reg  GEN_6;
  reg [31:0] GEN_14;
  reg [2:0] GEN_7;
  reg [31:0] GEN_15;
  reg [63:0] GEN_8;
  reg [63:0] GEN_16;
  FinishUnit finisher (
    .clk(finisher_clk),
    .reset(finisher_reset),
    .io_grant_ready(finisher_io_grant_ready),
    .io_grant_valid(finisher_io_grant_valid),
    .io_grant_bits_header_src(finisher_io_grant_bits_header_src),
    .io_grant_bits_header_dst(finisher_io_grant_bits_header_dst),
    .io_grant_bits_payload_addr_beat(finisher_io_grant_bits_payload_addr_beat),
    .io_grant_bits_payload_client_xact_id(finisher_io_grant_bits_payload_client_xact_id),
    .io_grant_bits_payload_manager_xact_id(finisher_io_grant_bits_payload_manager_xact_id),
    .io_grant_bits_payload_is_builtin_type(finisher_io_grant_bits_payload_is_builtin_type),
    .io_grant_bits_payload_g_type(finisher_io_grant_bits_payload_g_type),
    .io_grant_bits_payload_data(finisher_io_grant_bits_payload_data),
    .io_refill_ready(finisher_io_refill_ready),
    .io_refill_valid(finisher_io_refill_valid),
    .io_refill_bits_addr_beat(finisher_io_refill_bits_addr_beat),
    .io_refill_bits_client_xact_id(finisher_io_refill_bits_client_xact_id),
    .io_refill_bits_manager_xact_id(finisher_io_refill_bits_manager_xact_id),
    .io_refill_bits_is_builtin_type(finisher_io_refill_bits_is_builtin_type),
    .io_refill_bits_g_type(finisher_io_refill_bits_g_type),
    .io_refill_bits_data(finisher_io_refill_bits_data),
    .io_finish_ready(finisher_io_finish_ready),
    .io_finish_valid(finisher_io_finish_valid),
    .io_finish_bits_header_src(finisher_io_finish_bits_header_src),
    .io_finish_bits_header_dst(finisher_io_finish_bits_header_dst),
    .io_finish_bits_payload_manager_xact_id(finisher_io_finish_bits_payload_manager_xact_id),
    .io_ready(finisher_io_ready)
  );
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_network_acquire_valid = T_3774;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_probe_ready = 1'h0;
  assign io_network_release_valid = 1'h0;
  assign io_network_release_bits_header_src = GEN_1;
  assign io_network_release_bits_header_dst = GEN_2;
  assign io_network_release_bits_payload_addr_beat = GEN_3;
  assign io_network_release_bits_payload_addr_block = GEN_4;
  assign io_network_release_bits_payload_client_xact_id = GEN_5;
  assign io_network_release_bits_payload_voluntary = GEN_6;
  assign io_network_release_bits_payload_r_type = GEN_7;
  assign io_network_release_bits_payload_data = GEN_8;
  assign finisher_clk = clk;
  assign finisher_reset = reset;
  assign finisher_io_grant_valid = io_network_grant_valid;
  assign finisher_io_grant_bits_header_src = io_network_grant_bits_header_src;
  assign finisher_io_grant_bits_header_dst = io_network_grant_bits_header_dst;
  assign finisher_io_grant_bits_payload_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign finisher_io_grant_bits_payload_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign finisher_io_grant_bits_payload_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign finisher_io_grant_bits_payload_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign finisher_io_grant_bits_payload_g_type = io_network_grant_bits_payload_g_type;
  assign finisher_io_grant_bits_payload_data = io_network_grant_bits_payload_data;
  assign finisher_io_refill_ready = io_client_grant_ready;
  assign finisher_io_finish_ready = io_network_finish_ready;
  assign acq_with_header_ready = T_3775;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = {{1'd0}, 1'h1};
  assign acq_with_header_bits_header_dst = {{1'd0}, T_3773};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3765 = GEN_0 << 6;
  assign T_3767 = 32'h80000000 <= T_3765;
  assign T_3773 = T_3767 ? 1'h0 : 1'h1;
  assign T_3774 = acq_with_header_valid & finisher_io_ready;
  assign T_3775 = io_network_acquire_ready & finisher_io_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  GEN_1 = GEN_9[1:0];
  GEN_10 = {1{$random}};
  GEN_2 = GEN_10[1:0];
  GEN_11 = {1{$random}};
  GEN_3 = GEN_11[2:0];
  GEN_12 = {1{$random}};
  GEN_4 = GEN_12[25:0];
  GEN_13 = {1{$random}};
  GEN_5 = GEN_13[1:0];
  GEN_14 = {1{$random}};
  GEN_6 = GEN_14[0:0];
  GEN_15 = {1{$random}};
  GEN_7 = GEN_15[2:0];
  GEN_16 = {2{$random}};
  GEN_8 = GEN_16[63:0];
  end
`endif
endmodule
module ManagerTileLinkNetworkPort(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output [1:0] io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [11:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output  io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input  [1:0] io_manager_grant_bits_client_xact_id,
  input  [2:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input   io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input   io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output [1:0] io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output  io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [1:0] io_network_acquire_bits_header_src,
  input  [1:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input  [1:0] io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [11:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [1:0] io_network_grant_bits_header_src,
  output [1:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output [1:0] io_network_grant_bits_payload_client_xact_id,
  output [2:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [1:0] io_network_finish_bits_header_src,
  input  [1:0] io_network_finish_bits_header_dst,
  input  [2:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [1:0] io_network_probe_bits_header_src,
  output [1:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [1:0] io_network_release_bits_header_src,
  input  [1:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input  [1:0] io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6829_ready;
  wire  T_6829_valid;
  wire [1:0] T_6829_bits_header_src;
  wire [1:0] T_6829_bits_header_dst;
  wire [2:0] T_6829_bits_payload_addr_beat;
  wire [1:0] T_6829_bits_payload_client_xact_id;
  wire [2:0] T_6829_bits_payload_manager_xact_id;
  wire  T_6829_bits_payload_is_builtin_type;
  wire [3:0] T_6829_bits_payload_g_type;
  wire [63:0] T_6829_bits_payload_data;
  wire  T_6829_bits_payload_client_id;
  wire  T_7459_ready;
  wire  T_7459_valid;
  wire [1:0] T_7459_bits_header_src;
  wire [1:0] T_7459_bits_header_dst;
  wire [25:0] T_7459_bits_payload_addr_block;
  wire [1:0] T_7459_bits_payload_p_type;
  wire  T_7459_bits_payload_client_id;
  wire  T_7774_ready;
  wire  T_7774_valid;
  wire [25:0] T_7774_bits_addr_block;
  wire [1:0] T_7774_bits_client_xact_id;
  wire [2:0] T_7774_bits_addr_beat;
  wire  T_7774_bits_is_builtin_type;
  wire [2:0] T_7774_bits_a_type;
  wire [11:0] T_7774_bits_union;
  wire [63:0] T_7774_bits_data;
  wire  T_7902_ready;
  wire  T_7902_valid;
  wire [2:0] T_7902_bits_addr_beat;
  wire [25:0] T_7902_bits_addr_block;
  wire [1:0] T_7902_bits_client_xact_id;
  wire  T_7902_bits_voluntary;
  wire [2:0] T_7902_bits_r_type;
  wire [63:0] T_7902_bits_data;
  wire  T_8018_ready;
  wire  T_8018_valid;
  wire [2:0] T_8018_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_7774_valid;
  assign io_manager_acquire_bits_addr_block = T_7774_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_7774_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_7774_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_7774_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_7774_bits_a_type;
  assign io_manager_acquire_bits_union = T_7774_bits_union;
  assign io_manager_acquire_bits_data = T_7774_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[0];
  assign io_manager_grant_ready = T_6829_ready;
  assign io_manager_finish_valid = T_8018_valid;
  assign io_manager_finish_bits_manager_xact_id = T_8018_bits_manager_xact_id;
  assign io_manager_probe_ready = T_7459_ready;
  assign io_manager_release_valid = T_7902_valid;
  assign io_manager_release_bits_addr_beat = T_7902_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_7902_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_7902_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_7902_bits_voluntary;
  assign io_manager_release_bits_r_type = T_7902_bits_r_type;
  assign io_manager_release_bits_data = T_7902_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[0];
  assign io_network_acquire_ready = T_7774_ready;
  assign io_network_grant_valid = T_6829_valid;
  assign io_network_grant_bits_header_src = T_6829_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6829_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6829_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6829_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6829_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6829_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6829_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6829_bits_payload_data;
  assign io_network_finish_ready = T_8018_ready;
  assign io_network_probe_valid = T_7459_valid;
  assign io_network_probe_bits_header_src = T_7459_bits_header_src;
  assign io_network_probe_bits_header_dst = T_7459_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_7459_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_7459_bits_payload_p_type;
  assign io_network_release_ready = T_7902_ready;
  assign T_6829_ready = io_network_grant_ready;
  assign T_6829_valid = io_manager_grant_valid;
  assign T_6829_bits_header_src = {{1'd0}, 1'h0};
  assign T_6829_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6829_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6829_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6829_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6829_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6829_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6829_bits_payload_data = io_manager_grant_bits_data;
  assign T_6829_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_7459_ready = io_network_probe_ready;
  assign T_7459_valid = io_manager_probe_valid;
  assign T_7459_bits_header_src = {{1'd0}, 1'h0};
  assign T_7459_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_7459_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_7459_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_7459_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_7774_ready = io_manager_acquire_ready;
  assign T_7774_valid = io_network_acquire_valid;
  assign T_7774_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_7774_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_7774_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_7774_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_7774_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_7774_bits_union = io_network_acquire_bits_payload_union;
  assign T_7774_bits_data = io_network_acquire_bits_payload_data;
  assign T_7902_ready = io_manager_release_ready;
  assign T_7902_valid = io_network_release_valid;
  assign T_7902_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_7902_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_7902_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_7902_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_7902_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_7902_bits_data = io_network_release_bits_payload_data;
  assign T_8018_ready = io_manager_finish_ready;
  assign T_8018_valid = io_network_finish_valid;
  assign T_8018_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module TileLinkEnqueuer_2(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  assign io_client_acquire_ready = io_manager_acquire_ready;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_release_ready = io_manager_release_ready;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_release_valid = io_client_release_valid;
  assign io_manager_release_bits_header_src = io_client_release_bits_header_src;
  assign io_manager_release_bits_header_dst = io_client_release_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = io_client_release_bits_payload_data;
endmodule
module ManagerTileLinkNetworkPort_1(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output [1:0] io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [11:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output  io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input  [1:0] io_manager_grant_bits_client_xact_id,
  input  [2:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input   io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input   io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output [1:0] io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output  io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [1:0] io_network_acquire_bits_header_src,
  input  [1:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input  [1:0] io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [11:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [1:0] io_network_grant_bits_header_src,
  output [1:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output [1:0] io_network_grant_bits_payload_client_xact_id,
  output [2:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [1:0] io_network_finish_bits_header_src,
  input  [1:0] io_network_finish_bits_header_dst,
  input  [2:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [1:0] io_network_probe_bits_header_src,
  output [1:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [1:0] io_network_release_bits_header_src,
  input  [1:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input  [1:0] io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6829_ready;
  wire  T_6829_valid;
  wire [1:0] T_6829_bits_header_src;
  wire [1:0] T_6829_bits_header_dst;
  wire [2:0] T_6829_bits_payload_addr_beat;
  wire [1:0] T_6829_bits_payload_client_xact_id;
  wire [2:0] T_6829_bits_payload_manager_xact_id;
  wire  T_6829_bits_payload_is_builtin_type;
  wire [3:0] T_6829_bits_payload_g_type;
  wire [63:0] T_6829_bits_payload_data;
  wire  T_6829_bits_payload_client_id;
  wire  T_7459_ready;
  wire  T_7459_valid;
  wire [1:0] T_7459_bits_header_src;
  wire [1:0] T_7459_bits_header_dst;
  wire [25:0] T_7459_bits_payload_addr_block;
  wire [1:0] T_7459_bits_payload_p_type;
  wire  T_7459_bits_payload_client_id;
  wire  T_7774_ready;
  wire  T_7774_valid;
  wire [25:0] T_7774_bits_addr_block;
  wire [1:0] T_7774_bits_client_xact_id;
  wire [2:0] T_7774_bits_addr_beat;
  wire  T_7774_bits_is_builtin_type;
  wire [2:0] T_7774_bits_a_type;
  wire [11:0] T_7774_bits_union;
  wire [63:0] T_7774_bits_data;
  wire  T_7902_ready;
  wire  T_7902_valid;
  wire [2:0] T_7902_bits_addr_beat;
  wire [25:0] T_7902_bits_addr_block;
  wire [1:0] T_7902_bits_client_xact_id;
  wire  T_7902_bits_voluntary;
  wire [2:0] T_7902_bits_r_type;
  wire [63:0] T_7902_bits_data;
  wire  T_8018_ready;
  wire  T_8018_valid;
  wire [2:0] T_8018_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_7774_valid;
  assign io_manager_acquire_bits_addr_block = T_7774_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_7774_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_7774_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_7774_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_7774_bits_a_type;
  assign io_manager_acquire_bits_union = T_7774_bits_union;
  assign io_manager_acquire_bits_data = T_7774_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[0];
  assign io_manager_grant_ready = T_6829_ready;
  assign io_manager_finish_valid = T_8018_valid;
  assign io_manager_finish_bits_manager_xact_id = T_8018_bits_manager_xact_id;
  assign io_manager_probe_ready = T_7459_ready;
  assign io_manager_release_valid = T_7902_valid;
  assign io_manager_release_bits_addr_beat = T_7902_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_7902_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_7902_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_7902_bits_voluntary;
  assign io_manager_release_bits_r_type = T_7902_bits_r_type;
  assign io_manager_release_bits_data = T_7902_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[0];
  assign io_network_acquire_ready = T_7774_ready;
  assign io_network_grant_valid = T_6829_valid;
  assign io_network_grant_bits_header_src = T_6829_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6829_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6829_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6829_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6829_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6829_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6829_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6829_bits_payload_data;
  assign io_network_finish_ready = T_8018_ready;
  assign io_network_probe_valid = T_7459_valid;
  assign io_network_probe_bits_header_src = T_7459_bits_header_src;
  assign io_network_probe_bits_header_dst = T_7459_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_7459_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_7459_bits_payload_p_type;
  assign io_network_release_ready = T_7902_ready;
  assign T_6829_ready = io_network_grant_ready;
  assign T_6829_valid = io_manager_grant_valid;
  assign T_6829_bits_header_src = {{1'd0}, 1'h1};
  assign T_6829_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6829_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6829_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6829_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6829_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6829_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6829_bits_payload_data = io_manager_grant_bits_data;
  assign T_6829_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_7459_ready = io_network_probe_ready;
  assign T_7459_valid = io_manager_probe_valid;
  assign T_7459_bits_header_src = {{1'd0}, 1'h1};
  assign T_7459_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_7459_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_7459_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_7459_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_7774_ready = io_manager_acquire_ready;
  assign T_7774_valid = io_network_acquire_valid;
  assign T_7774_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_7774_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_7774_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_7774_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_7774_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_7774_bits_union = io_network_acquire_bits_payload_union;
  assign T_7774_bits_data = io_network_acquire_bits_payload_data;
  assign T_7902_ready = io_manager_release_ready;
  assign T_7902_valid = io_network_release_valid;
  assign T_7902_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_7902_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_7902_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_7902_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_7902_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_7902_bits_data = io_network_release_bits_payload_data;
  assign T_8018_ready = io_manager_finish_ready;
  assign T_8018_valid = io_network_finish_valid;
  assign T_8018_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module LockingRRArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [11:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [11:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [11:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [11:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_client_xact_id,
  output [2:0] io_out_bits_payload_addr_beat,
  output  io_out_bits_payload_is_builtin_type,
  output [2:0] io_out_bits_payload_a_type,
  output [11:0] io_out_bits_payload_union,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire [1:0] GEN_50;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_1;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire [1:0] GEN_2;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [25:0] GEN_3;
  wire [25:0] GEN_19;
  wire [25:0] GEN_20;
  wire [25:0] GEN_21;
  wire [1:0] GEN_4;
  wire [1:0] GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [2:0] GEN_5;
  wire [2:0] GEN_25;
  wire [2:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_6;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire [2:0] GEN_7;
  wire [2:0] GEN_31;
  wire [2:0] GEN_32;
  wire [2:0] GEN_33;
  wire [11:0] GEN_8;
  wire [11:0] GEN_34;
  wire [11:0] GEN_35;
  wire [11:0] GEN_36;
  wire [63:0] GEN_9;
  wire [63:0] GEN_37;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  reg [2:0] T_1236;
  reg [31:0] GEN_51;
  reg [1:0] T_1238;
  reg [31:0] GEN_52;
  wire [2:0] GEN_60;
  wire  T_1240;
  wire [2:0] T_1249_0;
  wire  T_1251;
  wire  T_1254;
  wire  T_1255;
  wire  T_1256;
  wire [2:0] GEN_61;
  wire [3:0] T_1260;
  wire [2:0] T_1261;
  wire [1:0] GEN_40;
  wire [2:0] GEN_41;
  wire [1:0] GEN_42;
  reg [1:0] lastGrant;
  reg [31:0] GEN_53;
  wire [1:0] GEN_43;
  wire  T_1266;
  wire  T_1268;
  wire  T_1270;
  wire  T_1272;
  wire  T_1273;
  wire  T_1274;
  wire  T_1277;
  wire  T_1278;
  wire  T_1279;
  wire  T_1280;
  wire  T_1281;
  wire  T_1285;
  wire  T_1287;
  wire  T_1289;
  wire  T_1291;
  wire  T_1293;
  wire  T_1295;
  wire  T_1299;
  wire  T_1300;
  wire  T_1301;
  wire  T_1302;
  wire  T_1303;
  wire [1:0] GEN_63;
  wire  T_1305;
  wire  T_1306;
  wire  T_1307;
  wire  T_1309;
  wire  T_1310;
  wire  T_1311;
  wire  T_1313;
  wire  T_1314;
  wire  T_1315;
  wire  T_1317;
  wire  T_1318;
  wire  T_1319;
  wire [1:0] GEN_44;
  wire [1:0] GEN_45;
  wire [1:0] GEN_46;
  wire [1:0] GEN_47;
  wire [1:0] GEN_48;
  wire [1:0] GEN_49;
  assign io_in_0_ready = T_1307;
  assign io_in_1_ready = T_1311;
  assign io_in_2_ready = T_1315;
  assign io_in_3_ready = T_1319;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_block = GEN_3;
  assign io_out_bits_payload_client_xact_id = GEN_4;
  assign io_out_bits_payload_addr_beat = GEN_5;
  assign io_out_bits_payload_is_builtin_type = GEN_6;
  assign io_out_bits_payload_a_type = GEN_7;
  assign io_out_bits_payload_union = GEN_8;
  assign io_out_bits_payload_data = GEN_9;
  assign io_chosen = GEN_42;
  assign choice = GEN_49;
  assign GEN_0 = GEN_12;
  assign GEN_50 = {{1'd0}, 1'h1};
  assign GEN_10 = GEN_50 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_valid : GEN_10;
  assign GEN_12 = 2'h3 == io_chosen ? io_in_3_valid : GEN_11;
  assign GEN_1 = GEN_15;
  assign GEN_13 = GEN_50 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_13;
  assign GEN_15 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_14;
  assign GEN_2 = GEN_18;
  assign GEN_16 = GEN_50 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_16;
  assign GEN_18 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_17;
  assign GEN_3 = GEN_21;
  assign GEN_19 = GEN_50 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_19;
  assign GEN_21 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_20;
  assign GEN_4 = GEN_24;
  assign GEN_22 = GEN_50 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_22;
  assign GEN_24 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_23;
  assign GEN_5 = GEN_27;
  assign GEN_25 = GEN_50 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_25;
  assign GEN_27 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_26;
  assign GEN_6 = GEN_30;
  assign GEN_28 = GEN_50 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_29 = 2'h2 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_28;
  assign GEN_30 = 2'h3 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_29;
  assign GEN_7 = GEN_33;
  assign GEN_31 = GEN_50 == io_chosen ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign GEN_32 = 2'h2 == io_chosen ? io_in_2_bits_payload_a_type : GEN_31;
  assign GEN_33 = 2'h3 == io_chosen ? io_in_3_bits_payload_a_type : GEN_32;
  assign GEN_8 = GEN_36;
  assign GEN_34 = GEN_50 == io_chosen ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign GEN_35 = 2'h2 == io_chosen ? io_in_2_bits_payload_union : GEN_34;
  assign GEN_36 = 2'h3 == io_chosen ? io_in_3_bits_payload_union : GEN_35;
  assign GEN_9 = GEN_39;
  assign GEN_37 = GEN_50 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_38 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_37;
  assign GEN_39 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_38;
  assign GEN_60 = {{2'd0}, 1'h0};
  assign T_1240 = T_1236 != GEN_60;
  assign T_1249_0 = 3'h3;
  assign T_1251 = T_1249_0 == io_out_bits_payload_a_type;
  assign T_1254 = io_out_bits_payload_is_builtin_type & T_1251;
  assign T_1255 = io_out_ready & io_out_valid;
  assign T_1256 = T_1255 & T_1254;
  assign GEN_61 = {{2'd0}, 1'h1};
  assign T_1260 = T_1236 + GEN_61;
  assign T_1261 = T_1260[2:0];
  assign GEN_40 = T_1256 ? io_chosen : T_1238;
  assign GEN_41 = T_1256 ? T_1261 : T_1236;
  assign GEN_42 = T_1240 ? T_1238 : choice;
  assign GEN_43 = T_1255 ? io_chosen : lastGrant;
  assign T_1266 = GEN_50 > lastGrant;
  assign T_1268 = 2'h2 > lastGrant;
  assign T_1270 = 2'h3 > lastGrant;
  assign T_1272 = io_in_1_valid & T_1266;
  assign T_1273 = io_in_2_valid & T_1268;
  assign T_1274 = io_in_3_valid & T_1270;
  assign T_1277 = T_1272 | T_1273;
  assign T_1278 = T_1277 | T_1274;
  assign T_1279 = T_1278 | io_in_0_valid;
  assign T_1280 = T_1279 | io_in_1_valid;
  assign T_1281 = T_1280 | io_in_2_valid;
  assign T_1285 = T_1272 == 1'h0;
  assign T_1287 = T_1277 == 1'h0;
  assign T_1289 = T_1278 == 1'h0;
  assign T_1291 = T_1279 == 1'h0;
  assign T_1293 = T_1280 == 1'h0;
  assign T_1295 = T_1281 == 1'h0;
  assign T_1299 = T_1266 | T_1291;
  assign T_1300 = T_1285 & T_1268;
  assign T_1301 = T_1300 | T_1293;
  assign T_1302 = T_1287 & T_1270;
  assign T_1303 = T_1302 | T_1295;
  assign GEN_63 = {{1'd0}, 1'h0};
  assign T_1305 = T_1238 == GEN_63;
  assign T_1306 = T_1240 ? T_1305 : T_1289;
  assign T_1307 = T_1306 & io_out_ready;
  assign T_1309 = T_1238 == GEN_50;
  assign T_1310 = T_1240 ? T_1309 : T_1299;
  assign T_1311 = T_1310 & io_out_ready;
  assign T_1313 = T_1238 == 2'h2;
  assign T_1314 = T_1240 ? T_1313 : T_1301;
  assign T_1315 = T_1314 & io_out_ready;
  assign T_1317 = T_1238 == 2'h3;
  assign T_1318 = T_1240 ? T_1317 : T_1303;
  assign T_1319 = T_1318 & io_out_ready;
  assign GEN_44 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_45 = io_in_1_valid ? {{1'd0}, 1'h1} : GEN_44;
  assign GEN_46 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_45;
  assign GEN_47 = T_1274 ? 2'h3 : GEN_46;
  assign GEN_48 = T_1273 ? 2'h2 : GEN_47;
  assign GEN_49 = T_1272 ? {{1'd0}, 1'h1} : GEN_48;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_51 = {1{$random}};
  T_1236 = GEN_51[2:0];
  GEN_52 = {1{$random}};
  T_1238 = GEN_52[1:0];
  GEN_53 = {1{$random}};
  lastGrant = GEN_53[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1236 <= 3'h0;
    end else begin
      if(T_1256) begin
        T_1236 <= T_1261;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1256) begin
        T_1238 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1255) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [11:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [11:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [11:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [11:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output  io_out_0_bits_payload_is_builtin_type,
  output [2:0] io_out_0_bits_payload_a_type,
  output [11:0] io_out_0_bits_payload_union,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output  io_out_1_bits_payload_is_builtin_type,
  output [2:0] io_out_1_bits_payload_a_type,
  output [11:0] io_out_1_bits_payload_union,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output  io_out_2_bits_payload_is_builtin_type,
  output [2:0] io_out_2_bits_payload_a_type,
  output [11:0] io_out_2_bits_payload_union,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output  io_out_3_bits_payload_is_builtin_type,
  output [2:0] io_out_3_bits_payload_a_type,
  output [11:0] io_out_3_bits_payload_union,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_0_bits_payload_a_type;
  wire [11:0] arb_io_in_0_bits_payload_union;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_1_bits_payload_a_type;
  wire [11:0] arb_io_in_1_bits_payload_union;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_2_bits_payload_a_type;
  wire [11:0] arb_io_in_2_bits_payload_union;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_3_bits_payload_a_type;
  wire [11:0] arb_io_in_3_bits_payload_union;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [2:0] arb_io_out_bits_payload_a_type;
  wire [11:0] arb_io_out_bits_payload_union;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire [1:0] GEN_4;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire [1:0] GEN_5;
  wire  T_1667;
  wire  T_1668;
  wire  T_1670;
  wire  T_1671;
  wire  T_1673;
  wire  T_1674;
  wire  T_1676;
  wire  T_1677;
  LockingRRArbiter arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(arb_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(arb_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(arb_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(arb_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(arb_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(arb_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(arb_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(arb_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_a_type(arb_io_out_bits_payload_a_type),
    .io_out_bits_payload_union(arb_io_out_bits_payload_union),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1668;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1671;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1674;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1677;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_3_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_a_type = io_in_0_bits_payload_a_type;
  assign arb_io_in_0_bits_payload_union = io_in_0_bits_payload_union;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_a_type = io_in_1_bits_payload_a_type;
  assign arb_io_in_1_bits_payload_union = io_in_1_bits_payload_union;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_a_type = io_in_2_bits_payload_a_type;
  assign arb_io_in_2_bits_payload_union = io_in_2_bits_payload_union;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_a_type = io_in_3_bits_payload_a_type;
  assign arb_io_in_3_bits_payload_union = io_in_3_bits_payload_union;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_4 = {{1'd0}, 1'h1};
  assign GEN_1 = GEN_4 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_5 = {{1'd0}, 1'h0};
  assign T_1667 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1668 = arb_io_out_valid & T_1667;
  assign T_1670 = arb_io_out_bits_header_dst == GEN_4;
  assign T_1671 = arb_io_out_valid & T_1670;
  assign T_1673 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1674 = arb_io_out_valid & T_1673;
  assign T_1676 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1677 = arb_io_out_valid & T_1676;
endmodule
module LockingRRArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_client_xact_id,
  output  io_out_bits_payload_voluntary,
  output [2:0] io_out_bits_payload_r_type,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire [1:0] GEN_46;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_1;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_2;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [2:0] GEN_3;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire [25:0] GEN_4;
  wire [25:0] GEN_21;
  wire [25:0] GEN_22;
  wire [25:0] GEN_23;
  wire [1:0] GEN_5;
  wire [1:0] GEN_24;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  wire  GEN_6;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire [2:0] GEN_7;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  wire [2:0] GEN_32;
  wire [63:0] GEN_8;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  reg [2:0] T_1202;
  reg [31:0] GEN_47;
  reg [1:0] T_1204;
  reg [31:0] GEN_48;
  wire [2:0] GEN_55;
  wire  T_1206;
  wire [2:0] T_1213_0;
  wire [2:0] T_1213_1;
  wire [2:0] T_1213_2;
  wire  T_1215;
  wire  T_1216;
  wire  T_1217;
  wire  T_1220;
  wire  T_1221;
  wire  T_1223;
  wire  T_1224;
  wire [2:0] GEN_56;
  wire [3:0] T_1228;
  wire [2:0] T_1229;
  wire [1:0] GEN_36;
  wire [2:0] GEN_37;
  wire [1:0] GEN_38;
  reg [1:0] lastGrant;
  reg [31:0] GEN_49;
  wire [1:0] GEN_39;
  wire  T_1234;
  wire  T_1236;
  wire  T_1238;
  wire  T_1240;
  wire  T_1241;
  wire  T_1242;
  wire  T_1245;
  wire  T_1246;
  wire  T_1247;
  wire  T_1248;
  wire  T_1249;
  wire  T_1253;
  wire  T_1255;
  wire  T_1257;
  wire  T_1259;
  wire  T_1261;
  wire  T_1263;
  wire  T_1267;
  wire  T_1268;
  wire  T_1269;
  wire  T_1270;
  wire  T_1271;
  wire [1:0] GEN_58;
  wire  T_1273;
  wire  T_1274;
  wire  T_1275;
  wire  T_1277;
  wire  T_1278;
  wire  T_1279;
  wire  T_1281;
  wire  T_1282;
  wire  T_1283;
  wire  T_1285;
  wire  T_1286;
  wire  T_1287;
  wire [1:0] GEN_40;
  wire [1:0] GEN_41;
  wire [1:0] GEN_42;
  wire [1:0] GEN_43;
  wire [1:0] GEN_44;
  wire [1:0] GEN_45;
  assign io_in_0_ready = T_1275;
  assign io_in_1_ready = T_1279;
  assign io_in_2_ready = T_1283;
  assign io_in_3_ready = T_1287;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_beat = GEN_3;
  assign io_out_bits_payload_addr_block = GEN_4;
  assign io_out_bits_payload_client_xact_id = GEN_5;
  assign io_out_bits_payload_voluntary = GEN_6;
  assign io_out_bits_payload_r_type = GEN_7;
  assign io_out_bits_payload_data = GEN_8;
  assign io_chosen = GEN_38;
  assign choice = GEN_45;
  assign GEN_0 = GEN_11;
  assign GEN_46 = {{1'd0}, 1'h1};
  assign GEN_9 = GEN_46 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 2'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_11 = 2'h3 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_1 = GEN_14;
  assign GEN_12 = GEN_46 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_12;
  assign GEN_14 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_13;
  assign GEN_2 = GEN_17;
  assign GEN_15 = GEN_46 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_15;
  assign GEN_17 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_16;
  assign GEN_3 = GEN_20;
  assign GEN_18 = GEN_46 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_18;
  assign GEN_20 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_19;
  assign GEN_4 = GEN_23;
  assign GEN_21 = GEN_46 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_21;
  assign GEN_23 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_22;
  assign GEN_5 = GEN_26;
  assign GEN_24 = GEN_46 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_24;
  assign GEN_26 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_25;
  assign GEN_6 = GEN_29;
  assign GEN_27 = GEN_46 == io_chosen ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_voluntary : GEN_27;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_bits_payload_voluntary : GEN_28;
  assign GEN_7 = GEN_32;
  assign GEN_30 = GEN_46 == io_chosen ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign GEN_31 = 2'h2 == io_chosen ? io_in_2_bits_payload_r_type : GEN_30;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_bits_payload_r_type : GEN_31;
  assign GEN_8 = GEN_35;
  assign GEN_33 = GEN_46 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_34 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_33;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_34;
  assign GEN_55 = {{2'd0}, 1'h0};
  assign T_1206 = T_1202 != GEN_55;
  assign T_1213_0 = 3'h0;
  assign T_1213_1 = 3'h1;
  assign T_1213_2 = 3'h2;
  assign T_1215 = T_1213_0 == io_out_bits_payload_r_type;
  assign T_1216 = T_1213_1 == io_out_bits_payload_r_type;
  assign T_1217 = T_1213_2 == io_out_bits_payload_r_type;
  assign T_1220 = T_1215 | T_1216;
  assign T_1221 = T_1220 | T_1217;
  assign T_1223 = io_out_ready & io_out_valid;
  assign T_1224 = T_1223 & T_1221;
  assign GEN_56 = {{2'd0}, 1'h1};
  assign T_1228 = T_1202 + GEN_56;
  assign T_1229 = T_1228[2:0];
  assign GEN_36 = T_1224 ? io_chosen : T_1204;
  assign GEN_37 = T_1224 ? T_1229 : T_1202;
  assign GEN_38 = T_1206 ? T_1204 : choice;
  assign GEN_39 = T_1223 ? io_chosen : lastGrant;
  assign T_1234 = GEN_46 > lastGrant;
  assign T_1236 = 2'h2 > lastGrant;
  assign T_1238 = 2'h3 > lastGrant;
  assign T_1240 = io_in_1_valid & T_1234;
  assign T_1241 = io_in_2_valid & T_1236;
  assign T_1242 = io_in_3_valid & T_1238;
  assign T_1245 = T_1240 | T_1241;
  assign T_1246 = T_1245 | T_1242;
  assign T_1247 = T_1246 | io_in_0_valid;
  assign T_1248 = T_1247 | io_in_1_valid;
  assign T_1249 = T_1248 | io_in_2_valid;
  assign T_1253 = T_1240 == 1'h0;
  assign T_1255 = T_1245 == 1'h0;
  assign T_1257 = T_1246 == 1'h0;
  assign T_1259 = T_1247 == 1'h0;
  assign T_1261 = T_1248 == 1'h0;
  assign T_1263 = T_1249 == 1'h0;
  assign T_1267 = T_1234 | T_1259;
  assign T_1268 = T_1253 & T_1236;
  assign T_1269 = T_1268 | T_1261;
  assign T_1270 = T_1255 & T_1238;
  assign T_1271 = T_1270 | T_1263;
  assign GEN_58 = {{1'd0}, 1'h0};
  assign T_1273 = T_1204 == GEN_58;
  assign T_1274 = T_1206 ? T_1273 : T_1257;
  assign T_1275 = T_1274 & io_out_ready;
  assign T_1277 = T_1204 == GEN_46;
  assign T_1278 = T_1206 ? T_1277 : T_1267;
  assign T_1279 = T_1278 & io_out_ready;
  assign T_1281 = T_1204 == 2'h2;
  assign T_1282 = T_1206 ? T_1281 : T_1269;
  assign T_1283 = T_1282 & io_out_ready;
  assign T_1285 = T_1204 == 2'h3;
  assign T_1286 = T_1206 ? T_1285 : T_1271;
  assign T_1287 = T_1286 & io_out_ready;
  assign GEN_40 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_41 = io_in_1_valid ? {{1'd0}, 1'h1} : GEN_40;
  assign GEN_42 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_41;
  assign GEN_43 = T_1242 ? 2'h3 : GEN_42;
  assign GEN_44 = T_1241 ? 2'h2 : GEN_43;
  assign GEN_45 = T_1240 ? {{1'd0}, 1'h1} : GEN_44;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_47 = {1{$random}};
  T_1202 = GEN_47[2:0];
  GEN_48 = {1{$random}};
  T_1204 = GEN_48[1:0];
  GEN_49 = {1{$random}};
  lastGrant = GEN_49[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1202 <= 3'h0;
    end else begin
      if(T_1224) begin
        T_1202 <= T_1229;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1224) begin
        T_1204 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1223) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output  io_out_0_bits_payload_voluntary,
  output [2:0] io_out_0_bits_payload_r_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output  io_out_1_bits_payload_voluntary,
  output [2:0] io_out_1_bits_payload_r_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output  io_out_2_bits_payload_voluntary,
  output [2:0] io_out_2_bits_payload_r_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output  io_out_3_bits_payload_voluntary,
  output [2:0] io_out_3_bits_payload_r_type,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire  arb_io_in_0_bits_payload_voluntary;
  wire [2:0] arb_io_in_0_bits_payload_r_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire  arb_io_in_1_bits_payload_voluntary;
  wire [2:0] arb_io_in_1_bits_payload_r_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire  arb_io_in_2_bits_payload_voluntary;
  wire [2:0] arb_io_in_2_bits_payload_r_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire  arb_io_in_3_bits_payload_voluntary;
  wire [2:0] arb_io_in_3_bits_payload_r_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire  arb_io_out_bits_payload_voluntary;
  wire [2:0] arb_io_out_bits_payload_r_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire [1:0] GEN_4;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire [1:0] GEN_5;
  wire  T_1621;
  wire  T_1622;
  wire  T_1624;
  wire  T_1625;
  wire  T_1627;
  wire  T_1628;
  wire  T_1630;
  wire  T_1631;
  LockingRRArbiter_1 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(arb_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(arb_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(arb_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(arb_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(arb_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(arb_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(arb_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(arb_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_voluntary(arb_io_out_bits_payload_voluntary),
    .io_out_bits_payload_r_type(arb_io_out_bits_payload_r_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1622;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_0_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1625;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_1_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1628;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_2_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1631;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_3_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_voluntary = io_in_0_bits_payload_voluntary;
  assign arb_io_in_0_bits_payload_r_type = io_in_0_bits_payload_r_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_voluntary = io_in_1_bits_payload_voluntary;
  assign arb_io_in_1_bits_payload_r_type = io_in_1_bits_payload_r_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_voluntary = io_in_2_bits_payload_voluntary;
  assign arb_io_in_2_bits_payload_r_type = io_in_2_bits_payload_r_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_voluntary = io_in_3_bits_payload_voluntary;
  assign arb_io_in_3_bits_payload_r_type = io_in_3_bits_payload_r_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_4 = {{1'd0}, 1'h1};
  assign GEN_1 = GEN_4 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_5 = {{1'd0}, 1'h0};
  assign T_1621 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1622 = arb_io_out_valid & T_1621;
  assign T_1624 = arb_io_out_bits_header_dst == GEN_4;
  assign T_1625 = arb_io_out_valid & T_1624;
  assign T_1627 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1628 = arb_io_out_valid & T_1627;
  assign T_1630 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1631 = arb_io_out_valid & T_1630;
endmodule
module LockingRRArbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_p_type,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire [1:0] GEN_27;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [1:0] GEN_1;
  wire [1:0] GEN_8;
  wire [1:0] GEN_9;
  wire [1:0] GEN_10;
  wire [1:0] GEN_2;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [25:0] GEN_3;
  wire [25:0] GEN_14;
  wire [25:0] GEN_15;
  wire [25:0] GEN_16;
  wire [1:0] GEN_4;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [1:0] GEN_19;
  wire  T_1066;
  reg [1:0] lastGrant;
  reg [31:0] GEN_28;
  wire [1:0] GEN_20;
  wire  T_1069;
  wire  T_1071;
  wire  T_1073;
  wire  T_1075;
  wire  T_1076;
  wire  T_1077;
  wire  T_1080;
  wire  T_1081;
  wire  T_1082;
  wire  T_1083;
  wire  T_1084;
  wire  T_1088;
  wire  T_1090;
  wire  T_1092;
  wire  T_1094;
  wire  T_1096;
  wire  T_1098;
  wire  T_1102;
  wire  T_1103;
  wire  T_1104;
  wire  T_1105;
  wire  T_1106;
  wire  T_1107;
  wire  T_1108;
  wire  T_1109;
  wire  T_1110;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  assign io_in_0_ready = T_1107;
  assign io_in_1_ready = T_1108;
  assign io_in_2_ready = T_1109;
  assign io_in_3_ready = T_1110;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_block = GEN_3;
  assign io_out_bits_payload_p_type = GEN_4;
  assign io_chosen = choice;
  assign choice = GEN_26;
  assign GEN_0 = GEN_7;
  assign GEN_27 = {{1'd0}, 1'h1};
  assign GEN_5 = GEN_27 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_6 = 2'h2 == io_chosen ? io_in_2_valid : GEN_5;
  assign GEN_7 = 2'h3 == io_chosen ? io_in_3_valid : GEN_6;
  assign GEN_1 = GEN_10;
  assign GEN_8 = GEN_27 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_9 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_8;
  assign GEN_10 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_9;
  assign GEN_2 = GEN_13;
  assign GEN_11 = GEN_27 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_12 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_11;
  assign GEN_13 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_12;
  assign GEN_3 = GEN_16;
  assign GEN_14 = GEN_27 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_14;
  assign GEN_16 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_15;
  assign GEN_4 = GEN_19;
  assign GEN_17 = GEN_27 == io_chosen ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_payload_p_type : GEN_17;
  assign GEN_19 = 2'h3 == io_chosen ? io_in_3_bits_payload_p_type : GEN_18;
  assign T_1066 = io_out_ready & io_out_valid;
  assign GEN_20 = T_1066 ? io_chosen : lastGrant;
  assign T_1069 = GEN_27 > lastGrant;
  assign T_1071 = 2'h2 > lastGrant;
  assign T_1073 = 2'h3 > lastGrant;
  assign T_1075 = io_in_1_valid & T_1069;
  assign T_1076 = io_in_2_valid & T_1071;
  assign T_1077 = io_in_3_valid & T_1073;
  assign T_1080 = T_1075 | T_1076;
  assign T_1081 = T_1080 | T_1077;
  assign T_1082 = T_1081 | io_in_0_valid;
  assign T_1083 = T_1082 | io_in_1_valid;
  assign T_1084 = T_1083 | io_in_2_valid;
  assign T_1088 = T_1075 == 1'h0;
  assign T_1090 = T_1080 == 1'h0;
  assign T_1092 = T_1081 == 1'h0;
  assign T_1094 = T_1082 == 1'h0;
  assign T_1096 = T_1083 == 1'h0;
  assign T_1098 = T_1084 == 1'h0;
  assign T_1102 = T_1069 | T_1094;
  assign T_1103 = T_1088 & T_1071;
  assign T_1104 = T_1103 | T_1096;
  assign T_1105 = T_1090 & T_1073;
  assign T_1106 = T_1105 | T_1098;
  assign T_1107 = T_1092 & io_out_ready;
  assign T_1108 = T_1102 & io_out_ready;
  assign T_1109 = T_1104 & io_out_ready;
  assign T_1110 = T_1106 & io_out_ready;
  assign GEN_21 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_22 = io_in_1_valid ? {{1'd0}, 1'h1} : GEN_21;
  assign GEN_23 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_22;
  assign GEN_24 = T_1077 ? 2'h3 : GEN_23;
  assign GEN_25 = T_1076 ? 2'h2 : GEN_24;
  assign GEN_26 = T_1075 ? {{1'd0}, 1'h1} : GEN_25;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_28 = {1{$random}};
  lastGrant = GEN_28[1:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_1066) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_p_type,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_p_type,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_p_type,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_p_type
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_p_type;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_p_type;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_p_type;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_p_type;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_p_type;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire [1:0] GEN_4;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire [1:0] GEN_5;
  wire  T_1437;
  wire  T_1438;
  wire  T_1440;
  wire  T_1441;
  wire  T_1443;
  wire  T_1444;
  wire  T_1446;
  wire  T_1447;
  LockingRRArbiter_2 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(arb_io_in_0_bits_payload_p_type),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(arb_io_in_1_bits_payload_p_type),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(arb_io_in_2_bits_payload_p_type),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(arb_io_in_3_bits_payload_p_type),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_p_type(arb_io_out_bits_payload_p_type),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1438;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_1_valid = T_1441;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_2_valid = T_1444;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_3_valid = T_1447;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_p_type = io_in_0_bits_payload_p_type;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_p_type = io_in_1_bits_payload_p_type;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_p_type = io_in_2_bits_payload_p_type;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_p_type = io_in_3_bits_payload_p_type;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_4 = {{1'd0}, 1'h1};
  assign GEN_1 = GEN_4 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_5 = {{1'd0}, 1'h0};
  assign T_1437 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1438 = arb_io_out_valid & T_1437;
  assign T_1440 = arb_io_out_bits_header_dst == GEN_4;
  assign T_1441 = arb_io_out_valid & T_1440;
  assign T_1443 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1444 = arb_io_out_valid & T_1443;
  assign T_1446 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1447 = arb_io_out_valid & T_1446;
endmodule
module LockingRRArbiter_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output [1:0] io_out_bits_payload_client_xact_id,
  output [2:0] io_out_bits_payload_manager_xact_id,
  output  io_out_bits_payload_is_builtin_type,
  output [3:0] io_out_bits_payload_g_type,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire [1:0] GEN_46;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_1;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_2;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [2:0] GEN_3;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire [1:0] GEN_4;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [1:0] GEN_23;
  wire [2:0] GEN_5;
  wire [2:0] GEN_24;
  wire [2:0] GEN_25;
  wire [2:0] GEN_26;
  wire  GEN_6;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire [3:0] GEN_7;
  wire [3:0] GEN_30;
  wire [3:0] GEN_31;
  wire [3:0] GEN_32;
  wire [63:0] GEN_8;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  reg [2:0] T_1202;
  reg [31:0] GEN_47;
  reg [1:0] T_1204;
  reg [31:0] GEN_48;
  wire [2:0] GEN_55;
  wire  T_1206;
  wire [2:0] T_1214_0;
  wire [3:0] GEN_56;
  wire  T_1216;
  wire [1:0] T_1224_0;
  wire [1:0] T_1224_1;
  wire [3:0] GEN_57;
  wire  T_1226;
  wire [3:0] GEN_58;
  wire  T_1227;
  wire  T_1230;
  wire  T_1231;
  wire  T_1233;
  wire  T_1234;
  wire [2:0] GEN_59;
  wire [3:0] T_1238;
  wire [2:0] T_1239;
  wire [1:0] GEN_36;
  wire [2:0] GEN_37;
  wire [1:0] GEN_38;
  reg [1:0] lastGrant;
  reg [31:0] GEN_49;
  wire [1:0] GEN_39;
  wire  T_1244;
  wire  T_1246;
  wire  T_1248;
  wire  T_1250;
  wire  T_1251;
  wire  T_1252;
  wire  T_1255;
  wire  T_1256;
  wire  T_1257;
  wire  T_1258;
  wire  T_1259;
  wire  T_1263;
  wire  T_1265;
  wire  T_1267;
  wire  T_1269;
  wire  T_1271;
  wire  T_1273;
  wire  T_1277;
  wire  T_1278;
  wire  T_1279;
  wire  T_1280;
  wire  T_1281;
  wire [1:0] GEN_61;
  wire  T_1283;
  wire  T_1284;
  wire  T_1285;
  wire  T_1287;
  wire  T_1288;
  wire  T_1289;
  wire  T_1291;
  wire  T_1292;
  wire  T_1293;
  wire  T_1295;
  wire  T_1296;
  wire  T_1297;
  wire [1:0] GEN_40;
  wire [1:0] GEN_41;
  wire [1:0] GEN_42;
  wire [1:0] GEN_43;
  wire [1:0] GEN_44;
  wire [1:0] GEN_45;
  assign io_in_0_ready = T_1285;
  assign io_in_1_ready = T_1289;
  assign io_in_2_ready = T_1293;
  assign io_in_3_ready = T_1297;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_beat = GEN_3;
  assign io_out_bits_payload_client_xact_id = GEN_4;
  assign io_out_bits_payload_manager_xact_id = GEN_5;
  assign io_out_bits_payload_is_builtin_type = GEN_6;
  assign io_out_bits_payload_g_type = GEN_7;
  assign io_out_bits_payload_data = GEN_8;
  assign io_chosen = GEN_38;
  assign choice = GEN_45;
  assign GEN_0 = GEN_11;
  assign GEN_46 = {{1'd0}, 1'h1};
  assign GEN_9 = GEN_46 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 2'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_11 = 2'h3 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_1 = GEN_14;
  assign GEN_12 = GEN_46 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_12;
  assign GEN_14 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_13;
  assign GEN_2 = GEN_17;
  assign GEN_15 = GEN_46 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_15;
  assign GEN_17 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_16;
  assign GEN_3 = GEN_20;
  assign GEN_18 = GEN_46 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_18;
  assign GEN_20 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_19;
  assign GEN_4 = GEN_23;
  assign GEN_21 = GEN_46 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_21;
  assign GEN_23 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_22;
  assign GEN_5 = GEN_26;
  assign GEN_24 = GEN_46 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_24;
  assign GEN_26 = 2'h3 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_25;
  assign GEN_6 = GEN_29;
  assign GEN_27 = GEN_46 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_27;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_28;
  assign GEN_7 = GEN_32;
  assign GEN_30 = GEN_46 == io_chosen ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign GEN_31 = 2'h2 == io_chosen ? io_in_2_bits_payload_g_type : GEN_30;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_bits_payload_g_type : GEN_31;
  assign GEN_8 = GEN_35;
  assign GEN_33 = GEN_46 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_34 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_33;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_34;
  assign GEN_55 = {{2'd0}, 1'h0};
  assign T_1206 = T_1202 != GEN_55;
  assign T_1214_0 = 3'h5;
  assign GEN_56 = {{1'd0}, T_1214_0};
  assign T_1216 = GEN_56 == io_out_bits_payload_g_type;
  assign T_1224_0 = 2'h0;
  assign T_1224_1 = 2'h1;
  assign GEN_57 = {{2'd0}, T_1224_0};
  assign T_1226 = GEN_57 == io_out_bits_payload_g_type;
  assign GEN_58 = {{2'd0}, T_1224_1};
  assign T_1227 = GEN_58 == io_out_bits_payload_g_type;
  assign T_1230 = T_1226 | T_1227;
  assign T_1231 = io_out_bits_payload_is_builtin_type ? T_1216 : T_1230;
  assign T_1233 = io_out_ready & io_out_valid;
  assign T_1234 = T_1233 & T_1231;
  assign GEN_59 = {{2'd0}, 1'h1};
  assign T_1238 = T_1202 + GEN_59;
  assign T_1239 = T_1238[2:0];
  assign GEN_36 = T_1234 ? io_chosen : T_1204;
  assign GEN_37 = T_1234 ? T_1239 : T_1202;
  assign GEN_38 = T_1206 ? T_1204 : choice;
  assign GEN_39 = T_1233 ? io_chosen : lastGrant;
  assign T_1244 = GEN_46 > lastGrant;
  assign T_1246 = 2'h2 > lastGrant;
  assign T_1248 = 2'h3 > lastGrant;
  assign T_1250 = io_in_1_valid & T_1244;
  assign T_1251 = io_in_2_valid & T_1246;
  assign T_1252 = io_in_3_valid & T_1248;
  assign T_1255 = T_1250 | T_1251;
  assign T_1256 = T_1255 | T_1252;
  assign T_1257 = T_1256 | io_in_0_valid;
  assign T_1258 = T_1257 | io_in_1_valid;
  assign T_1259 = T_1258 | io_in_2_valid;
  assign T_1263 = T_1250 == 1'h0;
  assign T_1265 = T_1255 == 1'h0;
  assign T_1267 = T_1256 == 1'h0;
  assign T_1269 = T_1257 == 1'h0;
  assign T_1271 = T_1258 == 1'h0;
  assign T_1273 = T_1259 == 1'h0;
  assign T_1277 = T_1244 | T_1269;
  assign T_1278 = T_1263 & T_1246;
  assign T_1279 = T_1278 | T_1271;
  assign T_1280 = T_1265 & T_1248;
  assign T_1281 = T_1280 | T_1273;
  assign GEN_61 = {{1'd0}, 1'h0};
  assign T_1283 = T_1204 == GEN_61;
  assign T_1284 = T_1206 ? T_1283 : T_1267;
  assign T_1285 = T_1284 & io_out_ready;
  assign T_1287 = T_1204 == GEN_46;
  assign T_1288 = T_1206 ? T_1287 : T_1277;
  assign T_1289 = T_1288 & io_out_ready;
  assign T_1291 = T_1204 == 2'h2;
  assign T_1292 = T_1206 ? T_1291 : T_1279;
  assign T_1293 = T_1292 & io_out_ready;
  assign T_1295 = T_1204 == 2'h3;
  assign T_1296 = T_1206 ? T_1295 : T_1281;
  assign T_1297 = T_1296 & io_out_ready;
  assign GEN_40 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_41 = io_in_1_valid ? {{1'd0}, 1'h1} : GEN_40;
  assign GEN_42 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_41;
  assign GEN_43 = T_1252 ? 2'h3 : GEN_42;
  assign GEN_44 = T_1251 ? 2'h2 : GEN_43;
  assign GEN_45 = T_1250 ? {{1'd0}, 1'h1} : GEN_44;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_47 = {1{$random}};
  T_1202 = GEN_47[2:0];
  GEN_48 = {1{$random}};
  T_1204 = GEN_48[1:0];
  GEN_49 = {1{$random}};
  lastGrant = GEN_49[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1202 <= 3'h0;
    end else begin
      if(T_1234) begin
        T_1202 <= T_1239;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1234) begin
        T_1204 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1233) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output [2:0] io_out_0_bits_payload_manager_xact_id,
  output  io_out_0_bits_payload_is_builtin_type,
  output [3:0] io_out_0_bits_payload_g_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output [2:0] io_out_1_bits_payload_manager_xact_id,
  output  io_out_1_bits_payload_is_builtin_type,
  output [3:0] io_out_1_bits_payload_g_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output [2:0] io_out_2_bits_payload_manager_xact_id,
  output  io_out_2_bits_payload_is_builtin_type,
  output [3:0] io_out_2_bits_payload_g_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output [2:0] io_out_3_bits_payload_manager_xact_id,
  output  io_out_3_bits_payload_is_builtin_type,
  output [3:0] io_out_3_bits_payload_g_type,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_0_bits_payload_g_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_1_bits_payload_g_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_2_bits_payload_g_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_3_bits_payload_g_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire [2:0] arb_io_out_bits_payload_manager_xact_id;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [3:0] arb_io_out_bits_payload_g_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire [1:0] GEN_4;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire [1:0] GEN_5;
  wire  T_1621;
  wire  T_1622;
  wire  T_1624;
  wire  T_1625;
  wire  T_1627;
  wire  T_1628;
  wire  T_1630;
  wire  T_1631;
  LockingRRArbiter_3 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(arb_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(arb_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(arb_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(arb_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_g_type(arb_io_out_bits_payload_g_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1622;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1625;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1628;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1631;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_g_type = io_in_0_bits_payload_g_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_g_type = io_in_1_bits_payload_g_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_g_type = io_in_2_bits_payload_g_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_g_type = io_in_3_bits_payload_g_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_4 = {{1'd0}, 1'h1};
  assign GEN_1 = GEN_4 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_5 = {{1'd0}, 1'h0};
  assign T_1621 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1622 = arb_io_out_valid & T_1621;
  assign T_1624 = arb_io_out_bits_header_dst == GEN_4;
  assign T_1625 = arb_io_out_valid & T_1624;
  assign T_1627 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1628 = arb_io_out_valid & T_1627;
  assign T_1630 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1631 = arb_io_out_valid & T_1630;
endmodule
module LockingRRArbiter_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_manager_xact_id,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire [1:0] GEN_23;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire [1:0] GEN_1;
  wire [1:0] GEN_7;
  wire [1:0] GEN_8;
  wire [1:0] GEN_9;
  wire [1:0] GEN_2;
  wire [1:0] GEN_10;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [2:0] GEN_3;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire  T_1032;
  reg [1:0] lastGrant;
  reg [31:0] GEN_24;
  wire [1:0] GEN_16;
  wire  T_1035;
  wire  T_1037;
  wire  T_1039;
  wire  T_1041;
  wire  T_1042;
  wire  T_1043;
  wire  T_1046;
  wire  T_1047;
  wire  T_1048;
  wire  T_1049;
  wire  T_1050;
  wire  T_1054;
  wire  T_1056;
  wire  T_1058;
  wire  T_1060;
  wire  T_1062;
  wire  T_1064;
  wire  T_1068;
  wire  T_1069;
  wire  T_1070;
  wire  T_1071;
  wire  T_1072;
  wire  T_1073;
  wire  T_1074;
  wire  T_1075;
  wire  T_1076;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [1:0] GEN_19;
  wire [1:0] GEN_20;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  assign io_in_0_ready = T_1073;
  assign io_in_1_ready = T_1074;
  assign io_in_2_ready = T_1075;
  assign io_in_3_ready = T_1076;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_manager_xact_id = GEN_3;
  assign io_chosen = choice;
  assign choice = GEN_22;
  assign GEN_0 = GEN_6;
  assign GEN_23 = {{1'd0}, 1'h1};
  assign GEN_4 = GEN_23 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_5 = 2'h2 == io_chosen ? io_in_2_valid : GEN_4;
  assign GEN_6 = 2'h3 == io_chosen ? io_in_3_valid : GEN_5;
  assign GEN_1 = GEN_9;
  assign GEN_7 = GEN_23 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_8 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_7;
  assign GEN_9 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_8;
  assign GEN_2 = GEN_12;
  assign GEN_10 = GEN_23 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_10;
  assign GEN_12 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_11;
  assign GEN_3 = GEN_15;
  assign GEN_13 = GEN_23 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_13;
  assign GEN_15 = 2'h3 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_14;
  assign T_1032 = io_out_ready & io_out_valid;
  assign GEN_16 = T_1032 ? io_chosen : lastGrant;
  assign T_1035 = GEN_23 > lastGrant;
  assign T_1037 = 2'h2 > lastGrant;
  assign T_1039 = 2'h3 > lastGrant;
  assign T_1041 = io_in_1_valid & T_1035;
  assign T_1042 = io_in_2_valid & T_1037;
  assign T_1043 = io_in_3_valid & T_1039;
  assign T_1046 = T_1041 | T_1042;
  assign T_1047 = T_1046 | T_1043;
  assign T_1048 = T_1047 | io_in_0_valid;
  assign T_1049 = T_1048 | io_in_1_valid;
  assign T_1050 = T_1049 | io_in_2_valid;
  assign T_1054 = T_1041 == 1'h0;
  assign T_1056 = T_1046 == 1'h0;
  assign T_1058 = T_1047 == 1'h0;
  assign T_1060 = T_1048 == 1'h0;
  assign T_1062 = T_1049 == 1'h0;
  assign T_1064 = T_1050 == 1'h0;
  assign T_1068 = T_1035 | T_1060;
  assign T_1069 = T_1054 & T_1037;
  assign T_1070 = T_1069 | T_1062;
  assign T_1071 = T_1056 & T_1039;
  assign T_1072 = T_1071 | T_1064;
  assign T_1073 = T_1058 & io_out_ready;
  assign T_1074 = T_1068 & io_out_ready;
  assign T_1075 = T_1070 & io_out_ready;
  assign T_1076 = T_1072 & io_out_ready;
  assign GEN_17 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_18 = io_in_1_valid ? {{1'd0}, 1'h1} : GEN_17;
  assign GEN_19 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_18;
  assign GEN_20 = T_1043 ? 2'h3 : GEN_19;
  assign GEN_21 = T_1042 ? 2'h2 : GEN_20;
  assign GEN_22 = T_1041 ? {{1'd0}, 1'h1} : GEN_21;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_24 = {1{$random}};
  lastGrant = GEN_24[1:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_1032) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_manager_xact_id,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_manager_xact_id,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_manager_xact_id,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_manager_xact_id
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_manager_xact_id;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire [1:0] GEN_4;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire [1:0] GEN_5;
  wire  T_1391;
  wire  T_1392;
  wire  T_1394;
  wire  T_1395;
  wire  T_1397;
  wire  T_1398;
  wire  T_1400;
  wire  T_1401;
  LockingRRArbiter_4 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1392;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_valid = T_1395;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_valid = T_1398;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_valid = T_1401;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_4 = {{1'd0}, 1'h1};
  assign GEN_1 = GEN_4 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_5 = {{1'd0}, 1'h0};
  assign T_1391 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1392 = arb_io_out_valid & T_1391;
  assign T_1394 = arb_io_out_bits_header_dst == GEN_4;
  assign T_1395 = arb_io_out_valid & T_1394;
  assign T_1397 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1398 = arb_io_out_valid & T_1397;
  assign T_1400 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1401 = arb_io_out_valid & T_1400;
endmodule
module PortedTileLinkCrossbar(
  input   clk,
  input   reset,
  output  io_clients_cached_0_acquire_ready,
  input   io_clients_cached_0_acquire_valid,
  input  [25:0] io_clients_cached_0_acquire_bits_addr_block,
  input  [1:0] io_clients_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_cached_0_acquire_bits_addr_beat,
  input   io_clients_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_cached_0_acquire_bits_a_type,
  input  [11:0] io_clients_cached_0_acquire_bits_union,
  input  [63:0] io_clients_cached_0_acquire_bits_data,
  input   io_clients_cached_0_probe_ready,
  output  io_clients_cached_0_probe_valid,
  output [25:0] io_clients_cached_0_probe_bits_addr_block,
  output [1:0] io_clients_cached_0_probe_bits_p_type,
  output  io_clients_cached_0_release_ready,
  input   io_clients_cached_0_release_valid,
  input  [2:0] io_clients_cached_0_release_bits_addr_beat,
  input  [25:0] io_clients_cached_0_release_bits_addr_block,
  input  [1:0] io_clients_cached_0_release_bits_client_xact_id,
  input   io_clients_cached_0_release_bits_voluntary,
  input  [2:0] io_clients_cached_0_release_bits_r_type,
  input  [63:0] io_clients_cached_0_release_bits_data,
  input   io_clients_cached_0_grant_ready,
  output  io_clients_cached_0_grant_valid,
  output [2:0] io_clients_cached_0_grant_bits_addr_beat,
  output [1:0] io_clients_cached_0_grant_bits_client_xact_id,
  output [2:0] io_clients_cached_0_grant_bits_manager_xact_id,
  output  io_clients_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_cached_0_grant_bits_g_type,
  output [63:0] io_clients_cached_0_grant_bits_data,
  output  io_clients_cached_0_grant_bits_manager_id,
  output  io_clients_cached_0_finish_ready,
  input   io_clients_cached_0_finish_valid,
  input  [2:0] io_clients_cached_0_finish_bits_manager_xact_id,
  input   io_clients_cached_0_finish_bits_manager_id,
  output  io_clients_uncached_0_acquire_ready,
  input   io_clients_uncached_0_acquire_valid,
  input  [25:0] io_clients_uncached_0_acquire_bits_addr_block,
  input  [1:0] io_clients_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_uncached_0_acquire_bits_addr_beat,
  input   io_clients_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_uncached_0_acquire_bits_a_type,
  input  [11:0] io_clients_uncached_0_acquire_bits_union,
  input  [63:0] io_clients_uncached_0_acquire_bits_data,
  input   io_clients_uncached_0_grant_ready,
  output  io_clients_uncached_0_grant_valid,
  output [2:0] io_clients_uncached_0_grant_bits_addr_beat,
  output [1:0] io_clients_uncached_0_grant_bits_client_xact_id,
  output [2:0] io_clients_uncached_0_grant_bits_manager_xact_id,
  output  io_clients_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_uncached_0_grant_bits_g_type,
  output [63:0] io_clients_uncached_0_grant_bits_data,
  input   io_managers_0_acquire_ready,
  output  io_managers_0_acquire_valid,
  output [25:0] io_managers_0_acquire_bits_addr_block,
  output [1:0] io_managers_0_acquire_bits_client_xact_id,
  output [2:0] io_managers_0_acquire_bits_addr_beat,
  output  io_managers_0_acquire_bits_is_builtin_type,
  output [2:0] io_managers_0_acquire_bits_a_type,
  output [11:0] io_managers_0_acquire_bits_union,
  output [63:0] io_managers_0_acquire_bits_data,
  output  io_managers_0_acquire_bits_client_id,
  output  io_managers_0_grant_ready,
  input   io_managers_0_grant_valid,
  input  [2:0] io_managers_0_grant_bits_addr_beat,
  input  [1:0] io_managers_0_grant_bits_client_xact_id,
  input  [2:0] io_managers_0_grant_bits_manager_xact_id,
  input   io_managers_0_grant_bits_is_builtin_type,
  input  [3:0] io_managers_0_grant_bits_g_type,
  input  [63:0] io_managers_0_grant_bits_data,
  input   io_managers_0_grant_bits_client_id,
  input   io_managers_0_finish_ready,
  output  io_managers_0_finish_valid,
  output [2:0] io_managers_0_finish_bits_manager_xact_id,
  output  io_managers_0_probe_ready,
  input   io_managers_0_probe_valid,
  input  [25:0] io_managers_0_probe_bits_addr_block,
  input  [1:0] io_managers_0_probe_bits_p_type,
  input   io_managers_0_probe_bits_client_id,
  input   io_managers_0_release_ready,
  output  io_managers_0_release_valid,
  output [2:0] io_managers_0_release_bits_addr_beat,
  output [25:0] io_managers_0_release_bits_addr_block,
  output [1:0] io_managers_0_release_bits_client_xact_id,
  output  io_managers_0_release_bits_voluntary,
  output [2:0] io_managers_0_release_bits_r_type,
  output [63:0] io_managers_0_release_bits_data,
  output  io_managers_0_release_bits_client_id,
  input   io_managers_1_acquire_ready,
  output  io_managers_1_acquire_valid,
  output [25:0] io_managers_1_acquire_bits_addr_block,
  output [1:0] io_managers_1_acquire_bits_client_xact_id,
  output [2:0] io_managers_1_acquire_bits_addr_beat,
  output  io_managers_1_acquire_bits_is_builtin_type,
  output [2:0] io_managers_1_acquire_bits_a_type,
  output [11:0] io_managers_1_acquire_bits_union,
  output [63:0] io_managers_1_acquire_bits_data,
  output  io_managers_1_acquire_bits_client_id,
  output  io_managers_1_grant_ready,
  input   io_managers_1_grant_valid,
  input  [2:0] io_managers_1_grant_bits_addr_beat,
  input  [1:0] io_managers_1_grant_bits_client_xact_id,
  input  [2:0] io_managers_1_grant_bits_manager_xact_id,
  input   io_managers_1_grant_bits_is_builtin_type,
  input  [3:0] io_managers_1_grant_bits_g_type,
  input  [63:0] io_managers_1_grant_bits_data,
  input   io_managers_1_grant_bits_client_id,
  input   io_managers_1_finish_ready,
  output  io_managers_1_finish_valid,
  output [2:0] io_managers_1_finish_bits_manager_xact_id,
  output  io_managers_1_probe_ready,
  input   io_managers_1_probe_valid,
  input  [25:0] io_managers_1_probe_bits_addr_block,
  input  [1:0] io_managers_1_probe_bits_p_type,
  input   io_managers_1_probe_bits_client_id,
  input   io_managers_1_release_ready,
  output  io_managers_1_release_valid,
  output [2:0] io_managers_1_release_bits_addr_beat,
  output [25:0] io_managers_1_release_bits_addr_block,
  output [1:0] io_managers_1_release_bits_client_xact_id,
  output  io_managers_1_release_bits_voluntary,
  output [2:0] io_managers_1_release_bits_r_type,
  output [63:0] io_managers_1_release_bits_data,
  output  io_managers_1_release_bits_client_id
);
  wire  TileLinkEnqueuer_4_clk;
  wire  TileLinkEnqueuer_4_reset;
  wire  TileLinkEnqueuer_4_io_client_acquire_ready;
  wire  TileLinkEnqueuer_4_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_client_grant_ready;
  wire  TileLinkEnqueuer_4_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_client_finish_ready;
  wire  TileLinkEnqueuer_4_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_client_probe_ready;
  wire  TileLinkEnqueuer_4_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_io_client_release_ready;
  wire  TileLinkEnqueuer_4_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_4_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_grant_ready;
  wire  TileLinkEnqueuer_4_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_finish_ready;
  wire  TileLinkEnqueuer_4_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_probe_ready;
  wire  TileLinkEnqueuer_4_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_io_manager_release_ready;
  wire  TileLinkEnqueuer_4_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_clk;
  wire  ClientTileLinkNetworkPort_1_reset;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_valid;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type;
  wire [11:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_union;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_probe_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_probe_valid;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  wire  ClientTileLinkNetworkPort_1_io_client_release_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_release_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_release_bits_r_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_release_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire [11:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_io_network_finish_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_finish_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_probe_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_probe_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire  ClientTileLinkNetworkPort_1_io_network_release_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_release_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_clk;
  wire  TileLinkEnqueuer_1_1_reset;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_1_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_1_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_1_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_1_1_io_client_release_ready;
  wire  TileLinkEnqueuer_1_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_1_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_clk;
  wire  ClientUncachedTileLinkNetworkPort_1_reset;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire [11:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_clk;
  wire  ManagerTileLinkNetworkPort_2_reset;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_finish_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_probe_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_clk;
  wire  TileLinkEnqueuer_2_1_reset;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_2_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_2_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_2_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_2_1_io_client_release_ready;
  wire  TileLinkEnqueuer_2_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_2_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_clk;
  wire  ManagerTileLinkNetworkPort_1_1_reset;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_probe_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_clk;
  wire  TileLinkEnqueuer_3_1_reset;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_3_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_3_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_3_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_3_1_io_client_release_ready;
  wire  TileLinkEnqueuer_3_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_3_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data;
  wire  acqNet_clk;
  wire  acqNet_reset;
  wire  acqNet_io_in_0_ready;
  wire  acqNet_io_in_0_valid;
  wire [1:0] acqNet_io_in_0_bits_header_src;
  wire [1:0] acqNet_io_in_0_bits_header_dst;
  wire [25:0] acqNet_io_in_0_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_0_bits_payload_addr_beat;
  wire  acqNet_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_0_bits_payload_a_type;
  wire [11:0] acqNet_io_in_0_bits_payload_union;
  wire [63:0] acqNet_io_in_0_bits_payload_data;
  wire  acqNet_io_in_1_ready;
  wire  acqNet_io_in_1_valid;
  wire [1:0] acqNet_io_in_1_bits_header_src;
  wire [1:0] acqNet_io_in_1_bits_header_dst;
  wire [25:0] acqNet_io_in_1_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_1_bits_payload_addr_beat;
  wire  acqNet_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_1_bits_payload_a_type;
  wire [11:0] acqNet_io_in_1_bits_payload_union;
  wire [63:0] acqNet_io_in_1_bits_payload_data;
  wire  acqNet_io_in_2_ready;
  wire  acqNet_io_in_2_valid;
  wire [1:0] acqNet_io_in_2_bits_header_src;
  wire [1:0] acqNet_io_in_2_bits_header_dst;
  wire [25:0] acqNet_io_in_2_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_2_bits_payload_addr_beat;
  wire  acqNet_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_2_bits_payload_a_type;
  wire [11:0] acqNet_io_in_2_bits_payload_union;
  wire [63:0] acqNet_io_in_2_bits_payload_data;
  wire  acqNet_io_in_3_ready;
  wire  acqNet_io_in_3_valid;
  wire [1:0] acqNet_io_in_3_bits_header_src;
  wire [1:0] acqNet_io_in_3_bits_header_dst;
  wire [25:0] acqNet_io_in_3_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_3_bits_payload_addr_beat;
  wire  acqNet_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_3_bits_payload_a_type;
  wire [11:0] acqNet_io_in_3_bits_payload_union;
  wire [63:0] acqNet_io_in_3_bits_payload_data;
  wire  acqNet_io_out_0_ready;
  wire  acqNet_io_out_0_valid;
  wire [1:0] acqNet_io_out_0_bits_header_src;
  wire [1:0] acqNet_io_out_0_bits_header_dst;
  wire [25:0] acqNet_io_out_0_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_0_bits_payload_addr_beat;
  wire  acqNet_io_out_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_0_bits_payload_a_type;
  wire [11:0] acqNet_io_out_0_bits_payload_union;
  wire [63:0] acqNet_io_out_0_bits_payload_data;
  wire  acqNet_io_out_1_ready;
  wire  acqNet_io_out_1_valid;
  wire [1:0] acqNet_io_out_1_bits_header_src;
  wire [1:0] acqNet_io_out_1_bits_header_dst;
  wire [25:0] acqNet_io_out_1_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_1_bits_payload_addr_beat;
  wire  acqNet_io_out_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_1_bits_payload_a_type;
  wire [11:0] acqNet_io_out_1_bits_payload_union;
  wire [63:0] acqNet_io_out_1_bits_payload_data;
  wire  acqNet_io_out_2_ready;
  wire  acqNet_io_out_2_valid;
  wire [1:0] acqNet_io_out_2_bits_header_src;
  wire [1:0] acqNet_io_out_2_bits_header_dst;
  wire [25:0] acqNet_io_out_2_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_2_bits_payload_addr_beat;
  wire  acqNet_io_out_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_2_bits_payload_a_type;
  wire [11:0] acqNet_io_out_2_bits_payload_union;
  wire [63:0] acqNet_io_out_2_bits_payload_data;
  wire  acqNet_io_out_3_ready;
  wire  acqNet_io_out_3_valid;
  wire [1:0] acqNet_io_out_3_bits_header_src;
  wire [1:0] acqNet_io_out_3_bits_header_dst;
  wire [25:0] acqNet_io_out_3_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_3_bits_payload_addr_beat;
  wire  acqNet_io_out_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_3_bits_payload_a_type;
  wire [11:0] acqNet_io_out_3_bits_payload_union;
  wire [63:0] acqNet_io_out_3_bits_payload_data;
  wire  relNet_clk;
  wire  relNet_reset;
  wire  relNet_io_in_0_ready;
  wire  relNet_io_in_0_valid;
  wire [1:0] relNet_io_in_0_bits_header_src;
  wire [1:0] relNet_io_in_0_bits_header_dst;
  wire [2:0] relNet_io_in_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_0_bits_payload_addr_block;
  wire [1:0] relNet_io_in_0_bits_payload_client_xact_id;
  wire  relNet_io_in_0_bits_payload_voluntary;
  wire [2:0] relNet_io_in_0_bits_payload_r_type;
  wire [63:0] relNet_io_in_0_bits_payload_data;
  wire  relNet_io_in_1_ready;
  wire  relNet_io_in_1_valid;
  wire [1:0] relNet_io_in_1_bits_header_src;
  wire [1:0] relNet_io_in_1_bits_header_dst;
  wire [2:0] relNet_io_in_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_1_bits_payload_addr_block;
  wire [1:0] relNet_io_in_1_bits_payload_client_xact_id;
  wire  relNet_io_in_1_bits_payload_voluntary;
  wire [2:0] relNet_io_in_1_bits_payload_r_type;
  wire [63:0] relNet_io_in_1_bits_payload_data;
  wire  relNet_io_in_2_ready;
  wire  relNet_io_in_2_valid;
  wire [1:0] relNet_io_in_2_bits_header_src;
  wire [1:0] relNet_io_in_2_bits_header_dst;
  wire [2:0] relNet_io_in_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_2_bits_payload_addr_block;
  wire [1:0] relNet_io_in_2_bits_payload_client_xact_id;
  wire  relNet_io_in_2_bits_payload_voluntary;
  wire [2:0] relNet_io_in_2_bits_payload_r_type;
  wire [63:0] relNet_io_in_2_bits_payload_data;
  wire  relNet_io_in_3_ready;
  wire  relNet_io_in_3_valid;
  wire [1:0] relNet_io_in_3_bits_header_src;
  wire [1:0] relNet_io_in_3_bits_header_dst;
  wire [2:0] relNet_io_in_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_3_bits_payload_addr_block;
  wire [1:0] relNet_io_in_3_bits_payload_client_xact_id;
  wire  relNet_io_in_3_bits_payload_voluntary;
  wire [2:0] relNet_io_in_3_bits_payload_r_type;
  wire [63:0] relNet_io_in_3_bits_payload_data;
  wire  relNet_io_out_0_ready;
  wire  relNet_io_out_0_valid;
  wire [1:0] relNet_io_out_0_bits_header_src;
  wire [1:0] relNet_io_out_0_bits_header_dst;
  wire [2:0] relNet_io_out_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_0_bits_payload_addr_block;
  wire [1:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire  relNet_io_out_0_bits_payload_voluntary;
  wire [2:0] relNet_io_out_0_bits_payload_r_type;
  wire [63:0] relNet_io_out_0_bits_payload_data;
  wire  relNet_io_out_1_ready;
  wire  relNet_io_out_1_valid;
  wire [1:0] relNet_io_out_1_bits_header_src;
  wire [1:0] relNet_io_out_1_bits_header_dst;
  wire [2:0] relNet_io_out_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_1_bits_payload_addr_block;
  wire [1:0] relNet_io_out_1_bits_payload_client_xact_id;
  wire  relNet_io_out_1_bits_payload_voluntary;
  wire [2:0] relNet_io_out_1_bits_payload_r_type;
  wire [63:0] relNet_io_out_1_bits_payload_data;
  wire  relNet_io_out_2_ready;
  wire  relNet_io_out_2_valid;
  wire [1:0] relNet_io_out_2_bits_header_src;
  wire [1:0] relNet_io_out_2_bits_header_dst;
  wire [2:0] relNet_io_out_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_2_bits_payload_addr_block;
  wire [1:0] relNet_io_out_2_bits_payload_client_xact_id;
  wire  relNet_io_out_2_bits_payload_voluntary;
  wire [2:0] relNet_io_out_2_bits_payload_r_type;
  wire [63:0] relNet_io_out_2_bits_payload_data;
  wire  relNet_io_out_3_ready;
  wire  relNet_io_out_3_valid;
  wire [1:0] relNet_io_out_3_bits_header_src;
  wire [1:0] relNet_io_out_3_bits_header_dst;
  wire [2:0] relNet_io_out_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_3_bits_payload_addr_block;
  wire [1:0] relNet_io_out_3_bits_payload_client_xact_id;
  wire  relNet_io_out_3_bits_payload_voluntary;
  wire [2:0] relNet_io_out_3_bits_payload_r_type;
  wire [63:0] relNet_io_out_3_bits_payload_data;
  wire  prbNet_clk;
  wire  prbNet_reset;
  wire  prbNet_io_in_0_ready;
  wire  prbNet_io_in_0_valid;
  wire [1:0] prbNet_io_in_0_bits_header_src;
  wire [1:0] prbNet_io_in_0_bits_header_dst;
  wire [25:0] prbNet_io_in_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_0_bits_payload_p_type;
  wire  prbNet_io_in_1_ready;
  wire  prbNet_io_in_1_valid;
  wire [1:0] prbNet_io_in_1_bits_header_src;
  wire [1:0] prbNet_io_in_1_bits_header_dst;
  wire [25:0] prbNet_io_in_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_1_bits_payload_p_type;
  wire  prbNet_io_in_2_ready;
  wire  prbNet_io_in_2_valid;
  wire [1:0] prbNet_io_in_2_bits_header_src;
  wire [1:0] prbNet_io_in_2_bits_header_dst;
  wire [25:0] prbNet_io_in_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_2_bits_payload_p_type;
  wire  prbNet_io_in_3_ready;
  wire  prbNet_io_in_3_valid;
  wire [1:0] prbNet_io_in_3_bits_header_src;
  wire [1:0] prbNet_io_in_3_bits_header_dst;
  wire [25:0] prbNet_io_in_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_3_bits_payload_p_type;
  wire  prbNet_io_out_0_ready;
  wire  prbNet_io_out_0_valid;
  wire [1:0] prbNet_io_out_0_bits_header_src;
  wire [1:0] prbNet_io_out_0_bits_header_dst;
  wire [25:0] prbNet_io_out_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_0_bits_payload_p_type;
  wire  prbNet_io_out_1_ready;
  wire  prbNet_io_out_1_valid;
  wire [1:0] prbNet_io_out_1_bits_header_src;
  wire [1:0] prbNet_io_out_1_bits_header_dst;
  wire [25:0] prbNet_io_out_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_1_bits_payload_p_type;
  wire  prbNet_io_out_2_ready;
  wire  prbNet_io_out_2_valid;
  wire [1:0] prbNet_io_out_2_bits_header_src;
  wire [1:0] prbNet_io_out_2_bits_header_dst;
  wire [25:0] prbNet_io_out_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_2_bits_payload_p_type;
  wire  prbNet_io_out_3_ready;
  wire  prbNet_io_out_3_valid;
  wire [1:0] prbNet_io_out_3_bits_header_src;
  wire [1:0] prbNet_io_out_3_bits_header_dst;
  wire [25:0] prbNet_io_out_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_3_bits_payload_p_type;
  wire  gntNet_clk;
  wire  gntNet_reset;
  wire  gntNet_io_in_0_ready;
  wire  gntNet_io_in_0_valid;
  wire [1:0] gntNet_io_in_0_bits_header_src;
  wire [1:0] gntNet_io_in_0_bits_header_dst;
  wire [2:0] gntNet_io_in_0_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_0_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_0_bits_payload_manager_xact_id;
  wire  gntNet_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_0_bits_payload_g_type;
  wire [63:0] gntNet_io_in_0_bits_payload_data;
  wire  gntNet_io_in_1_ready;
  wire  gntNet_io_in_1_valid;
  wire [1:0] gntNet_io_in_1_bits_header_src;
  wire [1:0] gntNet_io_in_1_bits_header_dst;
  wire [2:0] gntNet_io_in_1_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_1_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_1_bits_payload_manager_xact_id;
  wire  gntNet_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_1_bits_payload_g_type;
  wire [63:0] gntNet_io_in_1_bits_payload_data;
  wire  gntNet_io_in_2_ready;
  wire  gntNet_io_in_2_valid;
  wire [1:0] gntNet_io_in_2_bits_header_src;
  wire [1:0] gntNet_io_in_2_bits_header_dst;
  wire [2:0] gntNet_io_in_2_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_2_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_2_bits_payload_manager_xact_id;
  wire  gntNet_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_2_bits_payload_g_type;
  wire [63:0] gntNet_io_in_2_bits_payload_data;
  wire  gntNet_io_in_3_ready;
  wire  gntNet_io_in_3_valid;
  wire [1:0] gntNet_io_in_3_bits_header_src;
  wire [1:0] gntNet_io_in_3_bits_header_dst;
  wire [2:0] gntNet_io_in_3_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_3_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_3_bits_payload_manager_xact_id;
  wire  gntNet_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_3_bits_payload_g_type;
  wire [63:0] gntNet_io_in_3_bits_payload_data;
  wire  gntNet_io_out_0_ready;
  wire  gntNet_io_out_0_valid;
  wire [1:0] gntNet_io_out_0_bits_header_src;
  wire [1:0] gntNet_io_out_0_bits_header_dst;
  wire [2:0] gntNet_io_out_0_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_0_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_0_bits_payload_manager_xact_id;
  wire  gntNet_io_out_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_0_bits_payload_g_type;
  wire [63:0] gntNet_io_out_0_bits_payload_data;
  wire  gntNet_io_out_1_ready;
  wire  gntNet_io_out_1_valid;
  wire [1:0] gntNet_io_out_1_bits_header_src;
  wire [1:0] gntNet_io_out_1_bits_header_dst;
  wire [2:0] gntNet_io_out_1_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_1_bits_payload_manager_xact_id;
  wire  gntNet_io_out_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_1_bits_payload_g_type;
  wire [63:0] gntNet_io_out_1_bits_payload_data;
  wire  gntNet_io_out_2_ready;
  wire  gntNet_io_out_2_valid;
  wire [1:0] gntNet_io_out_2_bits_header_src;
  wire [1:0] gntNet_io_out_2_bits_header_dst;
  wire [2:0] gntNet_io_out_2_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_2_bits_payload_manager_xact_id;
  wire  gntNet_io_out_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_2_bits_payload_g_type;
  wire [63:0] gntNet_io_out_2_bits_payload_data;
  wire  gntNet_io_out_3_ready;
  wire  gntNet_io_out_3_valid;
  wire [1:0] gntNet_io_out_3_bits_header_src;
  wire [1:0] gntNet_io_out_3_bits_header_dst;
  wire [2:0] gntNet_io_out_3_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_3_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_3_bits_payload_manager_xact_id;
  wire  gntNet_io_out_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_3_bits_payload_g_type;
  wire [63:0] gntNet_io_out_3_bits_payload_data;
  wire  ackNet_clk;
  wire  ackNet_reset;
  wire  ackNet_io_in_0_ready;
  wire  ackNet_io_in_0_valid;
  wire [1:0] ackNet_io_in_0_bits_header_src;
  wire [1:0] ackNet_io_in_0_bits_header_dst;
  wire [2:0] ackNet_io_in_0_bits_payload_manager_xact_id;
  wire  ackNet_io_in_1_ready;
  wire  ackNet_io_in_1_valid;
  wire [1:0] ackNet_io_in_1_bits_header_src;
  wire [1:0] ackNet_io_in_1_bits_header_dst;
  wire [2:0] ackNet_io_in_1_bits_payload_manager_xact_id;
  wire  ackNet_io_in_2_ready;
  wire  ackNet_io_in_2_valid;
  wire [1:0] ackNet_io_in_2_bits_header_src;
  wire [1:0] ackNet_io_in_2_bits_header_dst;
  wire [2:0] ackNet_io_in_2_bits_payload_manager_xact_id;
  wire  ackNet_io_in_3_ready;
  wire  ackNet_io_in_3_valid;
  wire [1:0] ackNet_io_in_3_bits_header_src;
  wire [1:0] ackNet_io_in_3_bits_header_dst;
  wire [2:0] ackNet_io_in_3_bits_payload_manager_xact_id;
  wire  ackNet_io_out_0_ready;
  wire  ackNet_io_out_0_valid;
  wire [1:0] ackNet_io_out_0_bits_header_src;
  wire [1:0] ackNet_io_out_0_bits_header_dst;
  wire [2:0] ackNet_io_out_0_bits_payload_manager_xact_id;
  wire  ackNet_io_out_1_ready;
  wire  ackNet_io_out_1_valid;
  wire [1:0] ackNet_io_out_1_bits_header_src;
  wire [1:0] ackNet_io_out_1_bits_header_dst;
  wire [2:0] ackNet_io_out_1_bits_payload_manager_xact_id;
  wire  ackNet_io_out_2_ready;
  wire  ackNet_io_out_2_valid;
  wire [1:0] ackNet_io_out_2_bits_header_src;
  wire [1:0] ackNet_io_out_2_bits_header_dst;
  wire [2:0] ackNet_io_out_2_bits_payload_manager_xact_id;
  wire  ackNet_io_out_3_ready;
  wire  ackNet_io_out_3_valid;
  wire [1:0] ackNet_io_out_3_bits_header_src;
  wire [1:0] ackNet_io_out_3_bits_header_dst;
  wire [2:0] ackNet_io_out_3_bits_payload_manager_xact_id;
  wire  T_14149_ready;
  wire  T_14149_valid;
  wire [1:0] T_14149_bits_header_src;
  wire [1:0] T_14149_bits_header_dst;
  wire [25:0] T_14149_bits_payload_addr_block;
  wire [1:0] T_14149_bits_payload_client_xact_id;
  wire [2:0] T_14149_bits_payload_addr_beat;
  wire  T_14149_bits_payload_is_builtin_type;
  wire [2:0] T_14149_bits_payload_a_type;
  wire [11:0] T_14149_bits_payload_union;
  wire [63:0] T_14149_bits_payload_data;
  wire [2:0] T_14407;
  wire [1:0] T_14408;
  wire  T_14794_ready;
  wire  T_14794_valid;
  wire [1:0] T_14794_bits_header_src;
  wire [1:0] T_14794_bits_header_dst;
  wire [25:0] T_14794_bits_payload_addr_block;
  wire [1:0] T_14794_bits_payload_client_xact_id;
  wire [2:0] T_14794_bits_payload_addr_beat;
  wire  T_14794_bits_payload_is_builtin_type;
  wire [2:0] T_14794_bits_payload_a_type;
  wire [11:0] T_14794_bits_payload_union;
  wire [63:0] T_14794_bits_payload_data;
  wire [2:0] T_15052;
  wire [1:0] T_15053;
  wire  T_15163_ready;
  wire  T_15163_valid;
  wire [1:0] T_15163_bits_header_src;
  wire [1:0] T_15163_bits_header_dst;
  wire [25:0] T_15163_bits_payload_addr_block;
  wire [1:0] T_15163_bits_payload_client_xact_id;
  wire [2:0] T_15163_bits_payload_addr_beat;
  wire  T_15163_bits_payload_is_builtin_type;
  wire [2:0] T_15163_bits_payload_a_type;
  wire [11:0] T_15163_bits_payload_union;
  wire [63:0] T_15163_bits_payload_data;
  wire [2:0] T_15237;
  wire [1:0] T_15238;
  wire  T_15348_ready;
  wire  T_15348_valid;
  wire [1:0] T_15348_bits_header_src;
  wire [1:0] T_15348_bits_header_dst;
  wire [25:0] T_15348_bits_payload_addr_block;
  wire [1:0] T_15348_bits_payload_client_xact_id;
  wire [2:0] T_15348_bits_payload_addr_beat;
  wire  T_15348_bits_payload_is_builtin_type;
  wire [2:0] T_15348_bits_payload_a_type;
  wire [11:0] T_15348_bits_payload_union;
  wire [63:0] T_15348_bits_payload_data;
  wire [2:0] T_15422;
  wire [1:0] T_15423;
  wire  T_15806_ready;
  wire  T_15806_valid;
  wire [1:0] T_15806_bits_header_src;
  wire [1:0] T_15806_bits_header_dst;
  wire [2:0] T_15806_bits_payload_addr_beat;
  wire [25:0] T_15806_bits_payload_addr_block;
  wire [1:0] T_15806_bits_payload_client_xact_id;
  wire  T_15806_bits_payload_voluntary;
  wire [2:0] T_15806_bits_payload_r_type;
  wire [63:0] T_15806_bits_payload_data;
  wire [2:0] T_16062;
  wire [1:0] T_16063;
  wire  T_16446_ready;
  wire  T_16446_valid;
  wire [1:0] T_16446_bits_header_src;
  wire [1:0] T_16446_bits_header_dst;
  wire [2:0] T_16446_bits_payload_addr_beat;
  wire [25:0] T_16446_bits_payload_addr_block;
  wire [1:0] T_16446_bits_payload_client_xact_id;
  wire  T_16446_bits_payload_voluntary;
  wire [2:0] T_16446_bits_payload_r_type;
  wire [63:0] T_16446_bits_payload_data;
  wire [2:0] T_16702;
  wire [1:0] T_16703;
  wire  T_16810_ready;
  wire  T_16810_valid;
  wire [1:0] T_16810_bits_header_src;
  wire [1:0] T_16810_bits_header_dst;
  wire [2:0] T_16810_bits_payload_addr_beat;
  wire [25:0] T_16810_bits_payload_addr_block;
  wire [1:0] T_16810_bits_payload_client_xact_id;
  wire  T_16810_bits_payload_voluntary;
  wire [2:0] T_16810_bits_payload_r_type;
  wire [63:0] T_16810_bits_payload_data;
  wire [2:0] T_16882;
  wire [1:0] T_16883;
  wire  T_16990_ready;
  wire  T_16990_valid;
  wire [1:0] T_16990_bits_header_src;
  wire [1:0] T_16990_bits_header_dst;
  wire [2:0] T_16990_bits_payload_addr_beat;
  wire [25:0] T_16990_bits_payload_addr_block;
  wire [1:0] T_16990_bits_payload_client_xact_id;
  wire  T_16990_bits_payload_voluntary;
  wire [2:0] T_16990_bits_payload_r_type;
  wire [63:0] T_16990_bits_payload_data;
  wire [2:0] T_17062;
  wire [1:0] T_17063;
  wire  T_17158_ready;
  wire  T_17158_valid;
  wire [1:0] T_17158_bits_header_src;
  wire [1:0] T_17158_bits_header_dst;
  wire [25:0] T_17158_bits_payload_addr_block;
  wire [1:0] T_17158_bits_payload_p_type;
  wire [2:0] T_17222;
  wire [1:0] T_17223;
  wire  T_17318_ready;
  wire  T_17318_valid;
  wire [1:0] T_17318_bits_header_src;
  wire [1:0] T_17318_bits_header_dst;
  wire [25:0] T_17318_bits_payload_addr_block;
  wire [1:0] T_17318_bits_payload_p_type;
  wire [2:0] T_17382;
  wire [1:0] T_17383;
  wire  T_17754_ready;
  wire  T_17754_valid;
  wire [1:0] T_17754_bits_header_src;
  wire [1:0] T_17754_bits_header_dst;
  wire [25:0] T_17754_bits_payload_addr_block;
  wire [1:0] T_17754_bits_payload_p_type;
  wire [2:0] T_18002;
  wire [1:0] T_18003;
  wire  T_18374_ready;
  wire  T_18374_valid;
  wire [1:0] T_18374_bits_header_src;
  wire [1:0] T_18374_bits_header_dst;
  wire [25:0] T_18374_bits_payload_addr_block;
  wire [1:0] T_18374_bits_payload_p_type;
  wire [2:0] T_18622;
  wire [1:0] T_18623;
  wire  T_18730_ready;
  wire  T_18730_valid;
  wire [1:0] T_18730_bits_header_src;
  wire [1:0] T_18730_bits_header_dst;
  wire [2:0] T_18730_bits_payload_addr_beat;
  wire [1:0] T_18730_bits_payload_client_xact_id;
  wire [2:0] T_18730_bits_payload_manager_xact_id;
  wire  T_18730_bits_payload_is_builtin_type;
  wire [3:0] T_18730_bits_payload_g_type;
  wire [63:0] T_18730_bits_payload_data;
  wire [2:0] T_18802;
  wire [1:0] T_18803;
  wire  T_18910_ready;
  wire  T_18910_valid;
  wire [1:0] T_18910_bits_header_src;
  wire [1:0] T_18910_bits_header_dst;
  wire [2:0] T_18910_bits_payload_addr_beat;
  wire [1:0] T_18910_bits_payload_client_xact_id;
  wire [2:0] T_18910_bits_payload_manager_xact_id;
  wire  T_18910_bits_payload_is_builtin_type;
  wire [3:0] T_18910_bits_payload_g_type;
  wire [63:0] T_18910_bits_payload_data;
  wire [2:0] T_18982;
  wire [1:0] T_18983;
  wire  T_19366_ready;
  wire  T_19366_valid;
  wire [1:0] T_19366_bits_header_src;
  wire [1:0] T_19366_bits_header_dst;
  wire [2:0] T_19366_bits_payload_addr_beat;
  wire [1:0] T_19366_bits_payload_client_xact_id;
  wire [2:0] T_19366_bits_payload_manager_xact_id;
  wire  T_19366_bits_payload_is_builtin_type;
  wire [3:0] T_19366_bits_payload_g_type;
  wire [63:0] T_19366_bits_payload_data;
  wire [2:0] T_19622;
  wire [1:0] T_19623;
  wire  T_20006_ready;
  wire  T_20006_valid;
  wire [1:0] T_20006_bits_header_src;
  wire [1:0] T_20006_bits_header_dst;
  wire [2:0] T_20006_bits_payload_addr_beat;
  wire [1:0] T_20006_bits_payload_client_xact_id;
  wire [2:0] T_20006_bits_payload_manager_xact_id;
  wire  T_20006_bits_payload_is_builtin_type;
  wire [3:0] T_20006_bits_payload_g_type;
  wire [63:0] T_20006_bits_payload_data;
  wire [2:0] T_20262;
  wire [1:0] T_20263;
  wire  T_20631_ready;
  wire  T_20631_valid;
  wire [1:0] T_20631_bits_header_src;
  wire [1:0] T_20631_bits_header_dst;
  wire [2:0] T_20631_bits_payload_manager_xact_id;
  wire [2:0] T_20877;
  wire [1:0] T_20878;
  wire  T_21246_ready;
  wire  T_21246_valid;
  wire [1:0] T_21246_bits_header_src;
  wire [1:0] T_21246_bits_header_dst;
  wire [2:0] T_21246_bits_payload_manager_xact_id;
  wire [2:0] T_21492;
  wire [1:0] T_21493;
  wire  T_21585_ready;
  wire  T_21585_valid;
  wire [1:0] T_21585_bits_header_src;
  wire [1:0] T_21585_bits_header_dst;
  wire [2:0] T_21585_bits_payload_manager_xact_id;
  wire [2:0] T_21647;
  wire [1:0] T_21648;
  wire  T_21740_ready;
  wire  T_21740_valid;
  wire [1:0] T_21740_bits_header_src;
  wire [1:0] T_21740_bits_header_dst;
  wire [2:0] T_21740_bits_payload_manager_xact_id;
  wire [2:0] T_21802;
  wire [1:0] T_21803;
  reg [1:0] GEN_0;
  reg [31:0] GEN_64;
  reg [1:0] GEN_1;
  reg [31:0] GEN_65;
  reg [25:0] GEN_2;
  reg [31:0] GEN_66;
  reg [1:0] GEN_3;
  reg [31:0] GEN_67;
  reg [2:0] GEN_4;
  reg [31:0] GEN_68;
  reg  GEN_5;
  reg [31:0] GEN_69;
  reg [2:0] GEN_6;
  reg [31:0] GEN_70;
  reg [11:0] GEN_7;
  reg [31:0] GEN_71;
  reg [63:0] GEN_8;
  reg [63:0] GEN_72;
  reg [1:0] GEN_9;
  reg [31:0] GEN_73;
  reg [1:0] GEN_10;
  reg [31:0] GEN_74;
  reg [25:0] GEN_11;
  reg [31:0] GEN_75;
  reg [1:0] GEN_12;
  reg [31:0] GEN_76;
  reg [2:0] GEN_13;
  reg [31:0] GEN_77;
  reg  GEN_14;
  reg [31:0] GEN_78;
  reg [2:0] GEN_15;
  reg [31:0] GEN_79;
  reg [11:0] GEN_16;
  reg [31:0] GEN_80;
  reg [63:0] GEN_17;
  reg [63:0] GEN_81;
  reg [1:0] GEN_18;
  reg [31:0] GEN_82;
  reg [1:0] GEN_19;
  reg [31:0] GEN_83;
  reg [2:0] GEN_20;
  reg [31:0] GEN_84;
  reg [25:0] GEN_21;
  reg [31:0] GEN_85;
  reg [1:0] GEN_22;
  reg [31:0] GEN_86;
  reg  GEN_23;
  reg [31:0] GEN_87;
  reg [2:0] GEN_24;
  reg [31:0] GEN_88;
  reg [63:0] GEN_25;
  reg [63:0] GEN_89;
  reg [1:0] GEN_26;
  reg [31:0] GEN_90;
  reg [1:0] GEN_27;
  reg [31:0] GEN_91;
  reg [2:0] GEN_28;
  reg [31:0] GEN_92;
  reg [25:0] GEN_29;
  reg [31:0] GEN_93;
  reg [1:0] GEN_30;
  reg [31:0] GEN_94;
  reg  GEN_31;
  reg [31:0] GEN_95;
  reg [2:0] GEN_32;
  reg [31:0] GEN_96;
  reg [63:0] GEN_33;
  reg [63:0] GEN_97;
  reg [1:0] GEN_34;
  reg [31:0] GEN_98;
  reg [1:0] GEN_35;
  reg [31:0] GEN_99;
  reg [25:0] GEN_36;
  reg [31:0] GEN_100;
  reg [1:0] GEN_37;
  reg [31:0] GEN_101;
  reg [1:0] GEN_38;
  reg [31:0] GEN_102;
  reg [1:0] GEN_39;
  reg [31:0] GEN_103;
  reg [25:0] GEN_40;
  reg [31:0] GEN_104;
  reg [1:0] GEN_41;
  reg [31:0] GEN_105;
  reg [1:0] GEN_42;
  reg [31:0] GEN_106;
  reg [1:0] GEN_43;
  reg [31:0] GEN_107;
  reg [2:0] GEN_44;
  reg [31:0] GEN_108;
  reg [1:0] GEN_45;
  reg [31:0] GEN_109;
  reg [2:0] GEN_46;
  reg [31:0] GEN_110;
  reg  GEN_47;
  reg [31:0] GEN_111;
  reg [3:0] GEN_48;
  reg [31:0] GEN_112;
  reg [63:0] GEN_49;
  reg [63:0] GEN_113;
  reg [1:0] GEN_50;
  reg [31:0] GEN_114;
  reg [1:0] GEN_51;
  reg [31:0] GEN_115;
  reg [2:0] GEN_52;
  reg [31:0] GEN_116;
  reg [1:0] GEN_53;
  reg [31:0] GEN_117;
  reg [2:0] GEN_54;
  reg [31:0] GEN_118;
  reg  GEN_55;
  reg [31:0] GEN_119;
  reg [3:0] GEN_56;
  reg [31:0] GEN_120;
  reg [63:0] GEN_57;
  reg [63:0] GEN_121;
  reg [1:0] GEN_58;
  reg [31:0] GEN_122;
  reg [1:0] GEN_59;
  reg [31:0] GEN_123;
  reg [2:0] GEN_60;
  reg [31:0] GEN_124;
  reg [1:0] GEN_61;
  reg [31:0] GEN_125;
  reg [1:0] GEN_62;
  reg [31:0] GEN_126;
  reg [2:0] GEN_63;
  reg [31:0] GEN_127;
  TileLinkEnqueuer TileLinkEnqueuer_4 (
    .clk(TileLinkEnqueuer_4_clk),
    .reset(TileLinkEnqueuer_4_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_4_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_4_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_4_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_4_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_4_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_4_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_4_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_4_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_4_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_4_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_4_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_4_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_4_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_4_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_4_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_4_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_4_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_4_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_4_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_4_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_4_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_4_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_4_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_4_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_4_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_4_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_4_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_4_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_4_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_4_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_4_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_4_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_4_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_4_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_4_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_4_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_4_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_4_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_4_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_4_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_4_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_4_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_4_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_4_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_4_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_4_io_manager_release_bits_payload_data)
  );
  ClientTileLinkNetworkPort ClientTileLinkNetworkPort_1 (
    .clk(ClientTileLinkNetworkPort_1_clk),
    .reset(ClientTileLinkNetworkPort_1_reset),
    .io_client_acquire_ready(ClientTileLinkNetworkPort_1_io_client_acquire_ready),
    .io_client_acquire_valid(ClientTileLinkNetworkPort_1_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientTileLinkNetworkPort_1_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientTileLinkNetworkPort_1_io_client_acquire_bits_data),
    .io_client_probe_ready(ClientTileLinkNetworkPort_1_io_client_probe_ready),
    .io_client_probe_valid(ClientTileLinkNetworkPort_1_io_client_probe_valid),
    .io_client_probe_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block),
    .io_client_probe_bits_p_type(ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type),
    .io_client_release_ready(ClientTileLinkNetworkPort_1_io_client_release_ready),
    .io_client_release_valid(ClientTileLinkNetworkPort_1_io_client_release_valid),
    .io_client_release_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat),
    .io_client_release_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block),
    .io_client_release_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id),
    .io_client_release_bits_voluntary(ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary),
    .io_client_release_bits_r_type(ClientTileLinkNetworkPort_1_io_client_release_bits_r_type),
    .io_client_release_bits_data(ClientTileLinkNetworkPort_1_io_client_release_bits_data),
    .io_client_grant_ready(ClientTileLinkNetworkPort_1_io_client_grant_ready),
    .io_client_grant_valid(ClientTileLinkNetworkPort_1_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientTileLinkNetworkPort_1_io_client_grant_bits_data),
    .io_client_grant_bits_manager_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id),
    .io_client_finish_ready(ClientTileLinkNetworkPort_1_io_client_finish_ready),
    .io_client_finish_valid(ClientTileLinkNetworkPort_1_io_client_finish_valid),
    .io_client_finish_bits_manager_xact_id(ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id),
    .io_client_finish_bits_manager_id(ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id),
    .io_network_acquire_ready(ClientTileLinkNetworkPort_1_io_network_acquire_ready),
    .io_network_acquire_valid(ClientTileLinkNetworkPort_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientTileLinkNetworkPort_1_io_network_grant_ready),
    .io_network_grant_valid(ClientTileLinkNetworkPort_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientTileLinkNetworkPort_1_io_network_finish_ready),
    .io_network_finish_valid(ClientTileLinkNetworkPort_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientTileLinkNetworkPort_1_io_network_probe_ready),
    .io_network_probe_valid(ClientTileLinkNetworkPort_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientTileLinkNetworkPort_1_io_network_release_ready),
    .io_network_release_valid(ClientTileLinkNetworkPort_1_io_network_release_valid),
    .io_network_release_bits_header_src(ClientTileLinkNetworkPort_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_1_1 (
    .clk(TileLinkEnqueuer_1_1_clk),
    .reset(TileLinkEnqueuer_1_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_1_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_1_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_1_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_1_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_1_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_1_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_1_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_1_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_1_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_1_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_1_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_1_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_1_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_1_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_1_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_1_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_1_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_1_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_1_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_1_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_1_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_1_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_1_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_1_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_1_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_1_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_1_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data)
  );
  ClientUncachedTileLinkNetworkPort ClientUncachedTileLinkNetworkPort_1 (
    .clk(ClientUncachedTileLinkNetworkPort_1_clk),
    .reset(ClientUncachedTileLinkNetworkPort_1_reset),
    .io_client_acquire_ready(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready),
    .io_client_acquire_valid(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data),
    .io_client_grant_ready(ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready),
    .io_client_grant_valid(ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data),
    .io_network_acquire_ready(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready),
    .io_network_acquire_valid(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready),
    .io_network_grant_valid(ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready),
    .io_network_finish_valid(ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready),
    .io_network_probe_valid(ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientUncachedTileLinkNetworkPort_1_io_network_release_ready),
    .io_network_release_valid(ClientUncachedTileLinkNetworkPort_1_io_network_release_valid),
    .io_network_release_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort ManagerTileLinkNetworkPort_2 (
    .clk(ManagerTileLinkNetworkPort_2_clk),
    .reset(ManagerTileLinkNetworkPort_2_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_2_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_2_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_2_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_2_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_2_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_2_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_2_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_2_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_2_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_2_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_2_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_2_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_2_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_2_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_2_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_2_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_2_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_2_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_2_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_2_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_2_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_2_1 (
    .clk(TileLinkEnqueuer_2_1_clk),
    .reset(TileLinkEnqueuer_2_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_2_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_2_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_2_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_2_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_2_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_2_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_2_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_2_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_2_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_2_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_2_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_2_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_2_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_2_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_2_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_2_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_2_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_2_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_2_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_2_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_2_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_2_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_2_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_2_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_2_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_2_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_2_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort_1 ManagerTileLinkNetworkPort_1_1 (
    .clk(ManagerTileLinkNetworkPort_1_1_clk),
    .reset(ManagerTileLinkNetworkPort_1_1_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_1_1_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_1_1_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_1_1_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_1_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_1_1_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_1_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_1_1_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_1_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_1_1_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_1_1_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_3_1 (
    .clk(TileLinkEnqueuer_3_1_clk),
    .reset(TileLinkEnqueuer_3_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_3_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_3_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_3_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_3_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_3_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_3_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_3_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_3_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_3_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_3_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_3_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_3_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_3_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_3_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_3_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_3_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_3_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_3_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_3_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_3_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_3_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_3_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_3_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_3_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_3_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_3_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_3_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data)
  );
  BasicBus acqNet (
    .clk(acqNet_clk),
    .reset(acqNet_reset),
    .io_in_0_ready(acqNet_io_in_0_ready),
    .io_in_0_valid(acqNet_io_in_0_valid),
    .io_in_0_bits_header_src(acqNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(acqNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(acqNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(acqNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(acqNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(acqNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(acqNet_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(acqNet_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(acqNet_io_in_0_bits_payload_data),
    .io_in_1_ready(acqNet_io_in_1_ready),
    .io_in_1_valid(acqNet_io_in_1_valid),
    .io_in_1_bits_header_src(acqNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(acqNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(acqNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(acqNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(acqNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(acqNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(acqNet_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(acqNet_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(acqNet_io_in_1_bits_payload_data),
    .io_in_2_ready(acqNet_io_in_2_ready),
    .io_in_2_valid(acqNet_io_in_2_valid),
    .io_in_2_bits_header_src(acqNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(acqNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(acqNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(acqNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(acqNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(acqNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(acqNet_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(acqNet_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(acqNet_io_in_2_bits_payload_data),
    .io_in_3_ready(acqNet_io_in_3_ready),
    .io_in_3_valid(acqNet_io_in_3_valid),
    .io_in_3_bits_header_src(acqNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(acqNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(acqNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(acqNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(acqNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(acqNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(acqNet_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(acqNet_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(acqNet_io_in_3_bits_payload_data),
    .io_out_0_ready(acqNet_io_out_0_ready),
    .io_out_0_valid(acqNet_io_out_0_valid),
    .io_out_0_bits_header_src(acqNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(acqNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(acqNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(acqNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_addr_beat(acqNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_is_builtin_type(acqNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_a_type(acqNet_io_out_0_bits_payload_a_type),
    .io_out_0_bits_payload_union(acqNet_io_out_0_bits_payload_union),
    .io_out_0_bits_payload_data(acqNet_io_out_0_bits_payload_data),
    .io_out_1_ready(acqNet_io_out_1_ready),
    .io_out_1_valid(acqNet_io_out_1_valid),
    .io_out_1_bits_header_src(acqNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(acqNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(acqNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(acqNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_addr_beat(acqNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_is_builtin_type(acqNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_a_type(acqNet_io_out_1_bits_payload_a_type),
    .io_out_1_bits_payload_union(acqNet_io_out_1_bits_payload_union),
    .io_out_1_bits_payload_data(acqNet_io_out_1_bits_payload_data),
    .io_out_2_ready(acqNet_io_out_2_ready),
    .io_out_2_valid(acqNet_io_out_2_valid),
    .io_out_2_bits_header_src(acqNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(acqNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(acqNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(acqNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_addr_beat(acqNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_is_builtin_type(acqNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_a_type(acqNet_io_out_2_bits_payload_a_type),
    .io_out_2_bits_payload_union(acqNet_io_out_2_bits_payload_union),
    .io_out_2_bits_payload_data(acqNet_io_out_2_bits_payload_data),
    .io_out_3_ready(acqNet_io_out_3_ready),
    .io_out_3_valid(acqNet_io_out_3_valid),
    .io_out_3_bits_header_src(acqNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(acqNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(acqNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(acqNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_addr_beat(acqNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_is_builtin_type(acqNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_a_type(acqNet_io_out_3_bits_payload_a_type),
    .io_out_3_bits_payload_union(acqNet_io_out_3_bits_payload_union),
    .io_out_3_bits_payload_data(acqNet_io_out_3_bits_payload_data)
  );
  BasicBus_1 relNet (
    .clk(relNet_clk),
    .reset(relNet_reset),
    .io_in_0_ready(relNet_io_in_0_ready),
    .io_in_0_valid(relNet_io_in_0_valid),
    .io_in_0_bits_header_src(relNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(relNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(relNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(relNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(relNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(relNet_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(relNet_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(relNet_io_in_0_bits_payload_data),
    .io_in_1_ready(relNet_io_in_1_ready),
    .io_in_1_valid(relNet_io_in_1_valid),
    .io_in_1_bits_header_src(relNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(relNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(relNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(relNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(relNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(relNet_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(relNet_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(relNet_io_in_1_bits_payload_data),
    .io_in_2_ready(relNet_io_in_2_ready),
    .io_in_2_valid(relNet_io_in_2_valid),
    .io_in_2_bits_header_src(relNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(relNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(relNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(relNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(relNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(relNet_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(relNet_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(relNet_io_in_2_bits_payload_data),
    .io_in_3_ready(relNet_io_in_3_ready),
    .io_in_3_valid(relNet_io_in_3_valid),
    .io_in_3_bits_header_src(relNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(relNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(relNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(relNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(relNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(relNet_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(relNet_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(relNet_io_in_3_bits_payload_data),
    .io_out_0_ready(relNet_io_out_0_ready),
    .io_out_0_valid(relNet_io_out_0_valid),
    .io_out_0_bits_header_src(relNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(relNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(relNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_addr_block(relNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(relNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_voluntary(relNet_io_out_0_bits_payload_voluntary),
    .io_out_0_bits_payload_r_type(relNet_io_out_0_bits_payload_r_type),
    .io_out_0_bits_payload_data(relNet_io_out_0_bits_payload_data),
    .io_out_1_ready(relNet_io_out_1_ready),
    .io_out_1_valid(relNet_io_out_1_valid),
    .io_out_1_bits_header_src(relNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(relNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(relNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_addr_block(relNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(relNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_voluntary(relNet_io_out_1_bits_payload_voluntary),
    .io_out_1_bits_payload_r_type(relNet_io_out_1_bits_payload_r_type),
    .io_out_1_bits_payload_data(relNet_io_out_1_bits_payload_data),
    .io_out_2_ready(relNet_io_out_2_ready),
    .io_out_2_valid(relNet_io_out_2_valid),
    .io_out_2_bits_header_src(relNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(relNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(relNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_addr_block(relNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(relNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_voluntary(relNet_io_out_2_bits_payload_voluntary),
    .io_out_2_bits_payload_r_type(relNet_io_out_2_bits_payload_r_type),
    .io_out_2_bits_payload_data(relNet_io_out_2_bits_payload_data),
    .io_out_3_ready(relNet_io_out_3_ready),
    .io_out_3_valid(relNet_io_out_3_valid),
    .io_out_3_bits_header_src(relNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(relNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(relNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_addr_block(relNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(relNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_voluntary(relNet_io_out_3_bits_payload_voluntary),
    .io_out_3_bits_payload_r_type(relNet_io_out_3_bits_payload_r_type),
    .io_out_3_bits_payload_data(relNet_io_out_3_bits_payload_data)
  );
  BasicBus_2 prbNet (
    .clk(prbNet_clk),
    .reset(prbNet_reset),
    .io_in_0_ready(prbNet_io_in_0_ready),
    .io_in_0_valid(prbNet_io_in_0_valid),
    .io_in_0_bits_header_src(prbNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(prbNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(prbNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(prbNet_io_in_0_bits_payload_p_type),
    .io_in_1_ready(prbNet_io_in_1_ready),
    .io_in_1_valid(prbNet_io_in_1_valid),
    .io_in_1_bits_header_src(prbNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(prbNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(prbNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(prbNet_io_in_1_bits_payload_p_type),
    .io_in_2_ready(prbNet_io_in_2_ready),
    .io_in_2_valid(prbNet_io_in_2_valid),
    .io_in_2_bits_header_src(prbNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(prbNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(prbNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(prbNet_io_in_2_bits_payload_p_type),
    .io_in_3_ready(prbNet_io_in_3_ready),
    .io_in_3_valid(prbNet_io_in_3_valid),
    .io_in_3_bits_header_src(prbNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(prbNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(prbNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(prbNet_io_in_3_bits_payload_p_type),
    .io_out_0_ready(prbNet_io_out_0_ready),
    .io_out_0_valid(prbNet_io_out_0_valid),
    .io_out_0_bits_header_src(prbNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(prbNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(prbNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_p_type(prbNet_io_out_0_bits_payload_p_type),
    .io_out_1_ready(prbNet_io_out_1_ready),
    .io_out_1_valid(prbNet_io_out_1_valid),
    .io_out_1_bits_header_src(prbNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(prbNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(prbNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_p_type(prbNet_io_out_1_bits_payload_p_type),
    .io_out_2_ready(prbNet_io_out_2_ready),
    .io_out_2_valid(prbNet_io_out_2_valid),
    .io_out_2_bits_header_src(prbNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(prbNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(prbNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_p_type(prbNet_io_out_2_bits_payload_p_type),
    .io_out_3_ready(prbNet_io_out_3_ready),
    .io_out_3_valid(prbNet_io_out_3_valid),
    .io_out_3_bits_header_src(prbNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(prbNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(prbNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_p_type(prbNet_io_out_3_bits_payload_p_type)
  );
  BasicBus_3 gntNet (
    .clk(gntNet_clk),
    .reset(gntNet_reset),
    .io_in_0_ready(gntNet_io_in_0_ready),
    .io_in_0_valid(gntNet_io_in_0_valid),
    .io_in_0_bits_header_src(gntNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(gntNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(gntNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(gntNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(gntNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(gntNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(gntNet_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(gntNet_io_in_0_bits_payload_data),
    .io_in_1_ready(gntNet_io_in_1_ready),
    .io_in_1_valid(gntNet_io_in_1_valid),
    .io_in_1_bits_header_src(gntNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(gntNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(gntNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(gntNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(gntNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(gntNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(gntNet_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(gntNet_io_in_1_bits_payload_data),
    .io_in_2_ready(gntNet_io_in_2_ready),
    .io_in_2_valid(gntNet_io_in_2_valid),
    .io_in_2_bits_header_src(gntNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(gntNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(gntNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(gntNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(gntNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(gntNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(gntNet_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(gntNet_io_in_2_bits_payload_data),
    .io_in_3_ready(gntNet_io_in_3_ready),
    .io_in_3_valid(gntNet_io_in_3_valid),
    .io_in_3_bits_header_src(gntNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(gntNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(gntNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(gntNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(gntNet_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(gntNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(gntNet_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(gntNet_io_in_3_bits_payload_data),
    .io_out_0_ready(gntNet_io_out_0_ready),
    .io_out_0_valid(gntNet_io_out_0_valid),
    .io_out_0_bits_header_src(gntNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(gntNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(gntNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_client_xact_id(gntNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_manager_xact_id(gntNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_0_bits_payload_is_builtin_type(gntNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_g_type(gntNet_io_out_0_bits_payload_g_type),
    .io_out_0_bits_payload_data(gntNet_io_out_0_bits_payload_data),
    .io_out_1_ready(gntNet_io_out_1_ready),
    .io_out_1_valid(gntNet_io_out_1_valid),
    .io_out_1_bits_header_src(gntNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(gntNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(gntNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_client_xact_id(gntNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_manager_xact_id(gntNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_1_bits_payload_is_builtin_type(gntNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_g_type(gntNet_io_out_1_bits_payload_g_type),
    .io_out_1_bits_payload_data(gntNet_io_out_1_bits_payload_data),
    .io_out_2_ready(gntNet_io_out_2_ready),
    .io_out_2_valid(gntNet_io_out_2_valid),
    .io_out_2_bits_header_src(gntNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(gntNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(gntNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_client_xact_id(gntNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_manager_xact_id(gntNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_2_bits_payload_is_builtin_type(gntNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_g_type(gntNet_io_out_2_bits_payload_g_type),
    .io_out_2_bits_payload_data(gntNet_io_out_2_bits_payload_data),
    .io_out_3_ready(gntNet_io_out_3_ready),
    .io_out_3_valid(gntNet_io_out_3_valid),
    .io_out_3_bits_header_src(gntNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(gntNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(gntNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_client_xact_id(gntNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_manager_xact_id(gntNet_io_out_3_bits_payload_manager_xact_id),
    .io_out_3_bits_payload_is_builtin_type(gntNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_g_type(gntNet_io_out_3_bits_payload_g_type),
    .io_out_3_bits_payload_data(gntNet_io_out_3_bits_payload_data)
  );
  BasicBus_4 ackNet (
    .clk(ackNet_clk),
    .reset(ackNet_reset),
    .io_in_0_ready(ackNet_io_in_0_ready),
    .io_in_0_valid(ackNet_io_in_0_valid),
    .io_in_0_bits_header_src(ackNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(ackNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(ackNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(ackNet_io_in_1_ready),
    .io_in_1_valid(ackNet_io_in_1_valid),
    .io_in_1_bits_header_src(ackNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(ackNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(ackNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(ackNet_io_in_2_ready),
    .io_in_2_valid(ackNet_io_in_2_valid),
    .io_in_2_bits_header_src(ackNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(ackNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(ackNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(ackNet_io_in_3_ready),
    .io_in_3_valid(ackNet_io_in_3_valid),
    .io_in_3_bits_header_src(ackNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(ackNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(ackNet_io_in_3_bits_payload_manager_xact_id),
    .io_out_0_ready(ackNet_io_out_0_ready),
    .io_out_0_valid(ackNet_io_out_0_valid),
    .io_out_0_bits_header_src(ackNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(ackNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_manager_xact_id(ackNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_1_ready(ackNet_io_out_1_ready),
    .io_out_1_valid(ackNet_io_out_1_valid),
    .io_out_1_bits_header_src(ackNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(ackNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_manager_xact_id(ackNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_2_ready(ackNet_io_out_2_ready),
    .io_out_2_valid(ackNet_io_out_2_valid),
    .io_out_2_bits_header_src(ackNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(ackNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_manager_xact_id(ackNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_3_ready(ackNet_io_out_3_ready),
    .io_out_3_valid(ackNet_io_out_3_valid),
    .io_out_3_bits_header_src(ackNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(ackNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_manager_xact_id(ackNet_io_out_3_bits_payload_manager_xact_id)
  );
  assign io_clients_cached_0_acquire_ready = ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_cached_0_probe_valid = ClientTileLinkNetworkPort_1_io_client_probe_valid;
  assign io_clients_cached_0_probe_bits_addr_block = ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  assign io_clients_cached_0_probe_bits_p_type = ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  assign io_clients_cached_0_release_ready = ClientTileLinkNetworkPort_1_io_client_release_ready;
  assign io_clients_cached_0_grant_valid = ClientTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_cached_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_cached_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_cached_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_cached_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_cached_0_grant_bits_g_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_cached_0_grant_bits_data = ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_clients_cached_0_grant_bits_manager_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id;
  assign io_clients_cached_0_finish_ready = ClientTileLinkNetworkPort_1_io_client_finish_ready;
  assign io_clients_uncached_0_acquire_ready = ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_uncached_0_grant_valid = ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_uncached_0_grant_bits_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_uncached_0_grant_bits_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_uncached_0_grant_bits_manager_xact_id = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_uncached_0_grant_bits_is_builtin_type = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_uncached_0_grant_bits_g_type = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_uncached_0_grant_bits_data = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_2_io_manager_acquire_valid;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_2_io_manager_grant_ready;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_2_io_manager_finish_valid;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_2_io_manager_probe_ready;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_2_io_manager_release_valid;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_2_io_manager_release_bits_data;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id;
  assign io_managers_1_acquire_valid = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid;
  assign io_managers_1_acquire_bits_addr_block = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block;
  assign io_managers_1_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id;
  assign io_managers_1_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat;
  assign io_managers_1_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_1_acquire_bits_a_type = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type;
  assign io_managers_1_acquire_bits_union = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union;
  assign io_managers_1_acquire_bits_data = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data;
  assign io_managers_1_acquire_bits_client_id = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id;
  assign io_managers_1_grant_ready = ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready;
  assign io_managers_1_finish_valid = ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid;
  assign io_managers_1_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id;
  assign io_managers_1_probe_ready = ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready;
  assign io_managers_1_release_valid = ManagerTileLinkNetworkPort_1_1_io_manager_release_valid;
  assign io_managers_1_release_bits_addr_beat = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat;
  assign io_managers_1_release_bits_addr_block = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block;
  assign io_managers_1_release_bits_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id;
  assign io_managers_1_release_bits_voluntary = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary;
  assign io_managers_1_release_bits_r_type = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type;
  assign io_managers_1_release_bits_data = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data;
  assign io_managers_1_release_bits_client_id = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id;
  assign TileLinkEnqueuer_4_clk = clk;
  assign TileLinkEnqueuer_4_reset = reset;
  assign TileLinkEnqueuer_4_io_client_acquire_valid = ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_header_src = ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_union = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_data = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_4_io_client_grant_ready = ClientTileLinkNetworkPort_1_io_network_grant_ready;
  assign TileLinkEnqueuer_4_io_client_finish_valid = ClientTileLinkNetworkPort_1_io_network_finish_valid;
  assign TileLinkEnqueuer_4_io_client_finish_bits_header_src = ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_finish_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id = ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_io_client_probe_ready = ClientTileLinkNetworkPort_1_io_network_probe_ready;
  assign TileLinkEnqueuer_4_io_client_release_valid = ClientTileLinkNetworkPort_1_io_network_release_valid;
  assign TileLinkEnqueuer_4_io_client_release_bits_header_src = ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_release_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_r_type = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_data = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_4_io_manager_acquire_ready = T_15163_ready;
  assign TileLinkEnqueuer_4_io_manager_grant_valid = T_19366_valid;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_header_src = T_19366_bits_header_src;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_header_dst = T_19366_bits_header_dst;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat = T_19366_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id = T_19366_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id = T_19366_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type = T_19366_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type = T_19366_bits_payload_g_type;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_data = T_19366_bits_payload_data;
  assign TileLinkEnqueuer_4_io_manager_finish_ready = T_21585_ready;
  assign TileLinkEnqueuer_4_io_manager_probe_valid = T_17754_valid;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_header_src = T_17754_bits_header_src;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_header_dst = T_17754_bits_header_dst;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block = T_17754_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type = T_17754_bits_payload_p_type;
  assign TileLinkEnqueuer_4_io_manager_release_ready = T_16810_ready;
  assign ClientTileLinkNetworkPort_1_clk = clk;
  assign ClientTileLinkNetworkPort_1_reset = reset;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_valid = io_clients_cached_0_acquire_valid;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block = io_clients_cached_0_acquire_bits_addr_block;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id = io_clients_cached_0_acquire_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat = io_clients_cached_0_acquire_bits_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type = io_clients_cached_0_acquire_bits_is_builtin_type;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type = io_clients_cached_0_acquire_bits_a_type;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_union = io_clients_cached_0_acquire_bits_union;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_data = io_clients_cached_0_acquire_bits_data;
  assign ClientTileLinkNetworkPort_1_io_client_probe_ready = io_clients_cached_0_probe_ready;
  assign ClientTileLinkNetworkPort_1_io_client_release_valid = io_clients_cached_0_release_valid;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat = io_clients_cached_0_release_bits_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block = io_clients_cached_0_release_bits_addr_block;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id = io_clients_cached_0_release_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary = io_clients_cached_0_release_bits_voluntary;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_r_type = io_clients_cached_0_release_bits_r_type;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_data = io_clients_cached_0_release_bits_data;
  assign ClientTileLinkNetworkPort_1_io_client_grant_ready = io_clients_cached_0_grant_ready;
  assign ClientTileLinkNetworkPort_1_io_client_finish_valid = io_clients_cached_0_finish_valid;
  assign ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id = io_clients_cached_0_finish_bits_manager_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id = io_clients_cached_0_finish_bits_manager_id;
  assign ClientTileLinkNetworkPort_1_io_network_acquire_ready = TileLinkEnqueuer_4_io_client_acquire_ready;
  assign ClientTileLinkNetworkPort_1_io_network_grant_valid = TileLinkEnqueuer_4_io_client_grant_valid;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src = TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst = TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data = TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  assign ClientTileLinkNetworkPort_1_io_network_finish_ready = TileLinkEnqueuer_4_io_client_finish_ready;
  assign ClientTileLinkNetworkPort_1_io_network_probe_valid = TileLinkEnqueuer_4_io_client_probe_valid;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src = TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst = TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  assign ClientTileLinkNetworkPort_1_io_network_release_ready = TileLinkEnqueuer_4_io_client_release_ready;
  assign TileLinkEnqueuer_1_1_clk = clk;
  assign TileLinkEnqueuer_1_1_reset = reset;
  assign TileLinkEnqueuer_1_1_io_client_acquire_valid = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_client_grant_ready = ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready;
  assign TileLinkEnqueuer_1_1_io_client_finish_valid = ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_probe_ready = ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready;
  assign TileLinkEnqueuer_1_1_io_client_release_valid = ClientUncachedTileLinkNetworkPort_1_io_network_release_valid;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_data = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_manager_acquire_ready = T_15348_ready;
  assign TileLinkEnqueuer_1_1_io_manager_grant_valid = T_20006_valid;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src = T_20006_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst = T_20006_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat = T_20006_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id = T_20006_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id = T_20006_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type = T_20006_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type = T_20006_bits_payload_g_type;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data = T_20006_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_manager_finish_ready = T_21740_ready;
  assign TileLinkEnqueuer_1_1_io_manager_probe_valid = T_18374_valid;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src = T_18374_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst = T_18374_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block = T_18374_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type = T_18374_bits_payload_p_type;
  assign TileLinkEnqueuer_1_1_io_manager_release_ready = T_16990_ready;
  assign ClientUncachedTileLinkNetworkPort_1_clk = clk;
  assign ClientUncachedTileLinkNetworkPort_1_reset = reset;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid = io_clients_uncached_0_acquire_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block = io_clients_uncached_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id = io_clients_uncached_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat = io_clients_uncached_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type = io_clients_uncached_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type = io_clients_uncached_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union = io_clients_uncached_0_acquire_bits_union;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data = io_clients_uncached_0_acquire_bits_data;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready = io_clients_uncached_0_grant_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready = TileLinkEnqueuer_1_1_io_client_acquire_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid = TileLinkEnqueuer_1_1_io_client_grant_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src = TileLinkEnqueuer_1_1_io_client_grant_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst = TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready = TileLinkEnqueuer_1_1_io_client_finish_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid = TileLinkEnqueuer_1_1_io_client_probe_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src = TileLinkEnqueuer_1_1_io_client_probe_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst = TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_release_ready = TileLinkEnqueuer_1_1_io_client_release_ready;
  assign ManagerTileLinkNetworkPort_2_clk = clk;
  assign ManagerTileLinkNetworkPort_2_reset = reset;
  assign ManagerTileLinkNetworkPort_2_io_manager_acquire_ready = io_managers_0_acquire_ready;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_valid = io_managers_0_grant_valid;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat = io_managers_0_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id = io_managers_0_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id = io_managers_0_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type = io_managers_0_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type = io_managers_0_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data = io_managers_0_grant_bits_data;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id = io_managers_0_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_finish_ready = io_managers_0_finish_ready;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_valid = io_managers_0_probe_valid;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block = io_managers_0_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type = io_managers_0_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id = io_managers_0_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_release_ready = io_managers_0_release_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_valid = TileLinkEnqueuer_2_1_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src = TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_2_io_network_grant_ready = TileLinkEnqueuer_2_1_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_valid = TileLinkEnqueuer_2_1_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src = TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_probe_ready = TileLinkEnqueuer_2_1_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_release_valid = TileLinkEnqueuer_2_1_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src = TileLinkEnqueuer_2_1_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_2_1_clk = clk;
  assign TileLinkEnqueuer_2_1_reset = reset;
  assign TileLinkEnqueuer_2_1_io_client_acquire_valid = T_14149_valid;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src = T_14149_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst = T_14149_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block = T_14149_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id = T_14149_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat = T_14149_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type = T_14149_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type = T_14149_bits_payload_a_type;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union = T_14149_bits_payload_union;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data = T_14149_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_client_grant_ready = T_18730_ready;
  assign TileLinkEnqueuer_2_1_io_client_finish_valid = T_20631_valid;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_header_src = T_20631_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst = T_20631_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id = T_20631_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_probe_ready = T_17158_ready;
  assign TileLinkEnqueuer_2_1_io_client_release_valid = T_15806_valid;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_header_src = T_15806_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_header_dst = T_15806_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat = T_15806_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block = T_15806_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id = T_15806_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary = T_15806_bits_payload_voluntary;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type = T_15806_bits_payload_r_type;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_data = T_15806_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_manager_acquire_ready = ManagerTileLinkNetworkPort_2_io_network_acquire_ready;
  assign TileLinkEnqueuer_2_1_io_manager_grant_valid = ManagerTileLinkNetworkPort_2_io_network_grant_valid;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_manager_finish_ready = ManagerTileLinkNetworkPort_2_io_network_finish_ready;
  assign TileLinkEnqueuer_2_1_io_manager_probe_valid = ManagerTileLinkNetworkPort_2_io_network_probe_valid;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_2_1_io_manager_release_ready = ManagerTileLinkNetworkPort_2_io_network_release_ready;
  assign ManagerTileLinkNetworkPort_1_1_clk = clk;
  assign ManagerTileLinkNetworkPort_1_1_reset = reset;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready = io_managers_1_acquire_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid = io_managers_1_grant_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat = io_managers_1_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id = io_managers_1_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id = io_managers_1_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type = io_managers_1_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type = io_managers_1_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data = io_managers_1_grant_bits_data;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id = io_managers_1_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready = io_managers_1_finish_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid = io_managers_1_probe_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block = io_managers_1_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type = io_managers_1_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id = io_managers_1_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_release_ready = io_managers_1_release_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid = TileLinkEnqueuer_3_1_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src = TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_1_1_io_network_grant_ready = TileLinkEnqueuer_3_1_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_valid = TileLinkEnqueuer_3_1_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src = TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_probe_ready = TileLinkEnqueuer_3_1_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_valid = TileLinkEnqueuer_3_1_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src = TileLinkEnqueuer_3_1_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_3_1_clk = clk;
  assign TileLinkEnqueuer_3_1_reset = reset;
  assign TileLinkEnqueuer_3_1_io_client_acquire_valid = T_14794_valid;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src = T_14794_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst = T_14794_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block = T_14794_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id = T_14794_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat = T_14794_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type = T_14794_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type = T_14794_bits_payload_a_type;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union = T_14794_bits_payload_union;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data = T_14794_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_client_grant_ready = T_18910_ready;
  assign TileLinkEnqueuer_3_1_io_client_finish_valid = T_21246_valid;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_header_src = T_21246_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst = T_21246_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id = T_21246_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_probe_ready = T_17318_ready;
  assign TileLinkEnqueuer_3_1_io_client_release_valid = T_16446_valid;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_header_src = T_16446_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_header_dst = T_16446_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat = T_16446_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block = T_16446_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id = T_16446_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary = T_16446_bits_payload_voluntary;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type = T_16446_bits_payload_r_type;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_data = T_16446_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_manager_acquire_ready = ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready;
  assign TileLinkEnqueuer_3_1_io_manager_grant_valid = ManagerTileLinkNetworkPort_1_1_io_network_grant_valid;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_manager_finish_ready = ManagerTileLinkNetworkPort_1_1_io_network_finish_ready;
  assign TileLinkEnqueuer_3_1_io_manager_probe_valid = ManagerTileLinkNetworkPort_1_1_io_network_probe_valid;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_3_1_io_manager_release_ready = ManagerTileLinkNetworkPort_1_1_io_network_release_ready;
  assign acqNet_clk = clk;
  assign acqNet_reset = reset;
  assign acqNet_io_in_0_valid = 1'h0;
  assign acqNet_io_in_0_bits_header_src = GEN_0;
  assign acqNet_io_in_0_bits_header_dst = GEN_1;
  assign acqNet_io_in_0_bits_payload_addr_block = GEN_2;
  assign acqNet_io_in_0_bits_payload_client_xact_id = GEN_3;
  assign acqNet_io_in_0_bits_payload_addr_beat = GEN_4;
  assign acqNet_io_in_0_bits_payload_is_builtin_type = GEN_5;
  assign acqNet_io_in_0_bits_payload_a_type = GEN_6;
  assign acqNet_io_in_0_bits_payload_union = GEN_7;
  assign acqNet_io_in_0_bits_payload_data = GEN_8;
  assign acqNet_io_in_1_valid = 1'h0;
  assign acqNet_io_in_1_bits_header_src = GEN_9;
  assign acqNet_io_in_1_bits_header_dst = GEN_10;
  assign acqNet_io_in_1_bits_payload_addr_block = GEN_11;
  assign acqNet_io_in_1_bits_payload_client_xact_id = GEN_12;
  assign acqNet_io_in_1_bits_payload_addr_beat = GEN_13;
  assign acqNet_io_in_1_bits_payload_is_builtin_type = GEN_14;
  assign acqNet_io_in_1_bits_payload_a_type = GEN_15;
  assign acqNet_io_in_1_bits_payload_union = GEN_16;
  assign acqNet_io_in_1_bits_payload_data = GEN_17;
  assign acqNet_io_in_2_valid = T_15163_valid;
  assign acqNet_io_in_2_bits_header_src = T_15163_bits_header_src;
  assign acqNet_io_in_2_bits_header_dst = T_15163_bits_header_dst;
  assign acqNet_io_in_2_bits_payload_addr_block = T_15163_bits_payload_addr_block;
  assign acqNet_io_in_2_bits_payload_client_xact_id = T_15163_bits_payload_client_xact_id;
  assign acqNet_io_in_2_bits_payload_addr_beat = T_15163_bits_payload_addr_beat;
  assign acqNet_io_in_2_bits_payload_is_builtin_type = T_15163_bits_payload_is_builtin_type;
  assign acqNet_io_in_2_bits_payload_a_type = T_15163_bits_payload_a_type;
  assign acqNet_io_in_2_bits_payload_union = T_15163_bits_payload_union;
  assign acqNet_io_in_2_bits_payload_data = T_15163_bits_payload_data;
  assign acqNet_io_in_3_valid = T_15348_valid;
  assign acqNet_io_in_3_bits_header_src = T_15348_bits_header_src;
  assign acqNet_io_in_3_bits_header_dst = T_15348_bits_header_dst;
  assign acqNet_io_in_3_bits_payload_addr_block = T_15348_bits_payload_addr_block;
  assign acqNet_io_in_3_bits_payload_client_xact_id = T_15348_bits_payload_client_xact_id;
  assign acqNet_io_in_3_bits_payload_addr_beat = T_15348_bits_payload_addr_beat;
  assign acqNet_io_in_3_bits_payload_is_builtin_type = T_15348_bits_payload_is_builtin_type;
  assign acqNet_io_in_3_bits_payload_a_type = T_15348_bits_payload_a_type;
  assign acqNet_io_in_3_bits_payload_union = T_15348_bits_payload_union;
  assign acqNet_io_in_3_bits_payload_data = T_15348_bits_payload_data;
  assign acqNet_io_out_0_ready = T_14149_ready;
  assign acqNet_io_out_1_ready = T_14794_ready;
  assign acqNet_io_out_2_ready = 1'h0;
  assign acqNet_io_out_3_ready = 1'h0;
  assign relNet_clk = clk;
  assign relNet_reset = reset;
  assign relNet_io_in_0_valid = 1'h0;
  assign relNet_io_in_0_bits_header_src = GEN_18;
  assign relNet_io_in_0_bits_header_dst = GEN_19;
  assign relNet_io_in_0_bits_payload_addr_beat = GEN_20;
  assign relNet_io_in_0_bits_payload_addr_block = GEN_21;
  assign relNet_io_in_0_bits_payload_client_xact_id = GEN_22;
  assign relNet_io_in_0_bits_payload_voluntary = GEN_23;
  assign relNet_io_in_0_bits_payload_r_type = GEN_24;
  assign relNet_io_in_0_bits_payload_data = GEN_25;
  assign relNet_io_in_1_valid = 1'h0;
  assign relNet_io_in_1_bits_header_src = GEN_26;
  assign relNet_io_in_1_bits_header_dst = GEN_27;
  assign relNet_io_in_1_bits_payload_addr_beat = GEN_28;
  assign relNet_io_in_1_bits_payload_addr_block = GEN_29;
  assign relNet_io_in_1_bits_payload_client_xact_id = GEN_30;
  assign relNet_io_in_1_bits_payload_voluntary = GEN_31;
  assign relNet_io_in_1_bits_payload_r_type = GEN_32;
  assign relNet_io_in_1_bits_payload_data = GEN_33;
  assign relNet_io_in_2_valid = T_16810_valid;
  assign relNet_io_in_2_bits_header_src = T_16810_bits_header_src;
  assign relNet_io_in_2_bits_header_dst = T_16810_bits_header_dst;
  assign relNet_io_in_2_bits_payload_addr_beat = T_16810_bits_payload_addr_beat;
  assign relNet_io_in_2_bits_payload_addr_block = T_16810_bits_payload_addr_block;
  assign relNet_io_in_2_bits_payload_client_xact_id = T_16810_bits_payload_client_xact_id;
  assign relNet_io_in_2_bits_payload_voluntary = T_16810_bits_payload_voluntary;
  assign relNet_io_in_2_bits_payload_r_type = T_16810_bits_payload_r_type;
  assign relNet_io_in_2_bits_payload_data = T_16810_bits_payload_data;
  assign relNet_io_in_3_valid = T_16990_valid;
  assign relNet_io_in_3_bits_header_src = T_16990_bits_header_src;
  assign relNet_io_in_3_bits_header_dst = T_16990_bits_header_dst;
  assign relNet_io_in_3_bits_payload_addr_beat = T_16990_bits_payload_addr_beat;
  assign relNet_io_in_3_bits_payload_addr_block = T_16990_bits_payload_addr_block;
  assign relNet_io_in_3_bits_payload_client_xact_id = T_16990_bits_payload_client_xact_id;
  assign relNet_io_in_3_bits_payload_voluntary = T_16990_bits_payload_voluntary;
  assign relNet_io_in_3_bits_payload_r_type = T_16990_bits_payload_r_type;
  assign relNet_io_in_3_bits_payload_data = T_16990_bits_payload_data;
  assign relNet_io_out_0_ready = T_15806_ready;
  assign relNet_io_out_1_ready = T_16446_ready;
  assign relNet_io_out_2_ready = 1'h0;
  assign relNet_io_out_3_ready = 1'h0;
  assign prbNet_clk = clk;
  assign prbNet_reset = reset;
  assign prbNet_io_in_0_valid = T_17158_valid;
  assign prbNet_io_in_0_bits_header_src = T_17158_bits_header_src;
  assign prbNet_io_in_0_bits_header_dst = T_17158_bits_header_dst;
  assign prbNet_io_in_0_bits_payload_addr_block = T_17158_bits_payload_addr_block;
  assign prbNet_io_in_0_bits_payload_p_type = T_17158_bits_payload_p_type;
  assign prbNet_io_in_1_valid = T_17318_valid;
  assign prbNet_io_in_1_bits_header_src = T_17318_bits_header_src;
  assign prbNet_io_in_1_bits_header_dst = T_17318_bits_header_dst;
  assign prbNet_io_in_1_bits_payload_addr_block = T_17318_bits_payload_addr_block;
  assign prbNet_io_in_1_bits_payload_p_type = T_17318_bits_payload_p_type;
  assign prbNet_io_in_2_valid = 1'h0;
  assign prbNet_io_in_2_bits_header_src = GEN_34;
  assign prbNet_io_in_2_bits_header_dst = GEN_35;
  assign prbNet_io_in_2_bits_payload_addr_block = GEN_36;
  assign prbNet_io_in_2_bits_payload_p_type = GEN_37;
  assign prbNet_io_in_3_valid = 1'h0;
  assign prbNet_io_in_3_bits_header_src = GEN_38;
  assign prbNet_io_in_3_bits_header_dst = GEN_39;
  assign prbNet_io_in_3_bits_payload_addr_block = GEN_40;
  assign prbNet_io_in_3_bits_payload_p_type = GEN_41;
  assign prbNet_io_out_0_ready = 1'h0;
  assign prbNet_io_out_1_ready = 1'h0;
  assign prbNet_io_out_2_ready = T_17754_ready;
  assign prbNet_io_out_3_ready = T_18374_ready;
  assign gntNet_clk = clk;
  assign gntNet_reset = reset;
  assign gntNet_io_in_0_valid = T_18730_valid;
  assign gntNet_io_in_0_bits_header_src = T_18730_bits_header_src;
  assign gntNet_io_in_0_bits_header_dst = T_18730_bits_header_dst;
  assign gntNet_io_in_0_bits_payload_addr_beat = T_18730_bits_payload_addr_beat;
  assign gntNet_io_in_0_bits_payload_client_xact_id = T_18730_bits_payload_client_xact_id;
  assign gntNet_io_in_0_bits_payload_manager_xact_id = T_18730_bits_payload_manager_xact_id;
  assign gntNet_io_in_0_bits_payload_is_builtin_type = T_18730_bits_payload_is_builtin_type;
  assign gntNet_io_in_0_bits_payload_g_type = T_18730_bits_payload_g_type;
  assign gntNet_io_in_0_bits_payload_data = T_18730_bits_payload_data;
  assign gntNet_io_in_1_valid = T_18910_valid;
  assign gntNet_io_in_1_bits_header_src = T_18910_bits_header_src;
  assign gntNet_io_in_1_bits_header_dst = T_18910_bits_header_dst;
  assign gntNet_io_in_1_bits_payload_addr_beat = T_18910_bits_payload_addr_beat;
  assign gntNet_io_in_1_bits_payload_client_xact_id = T_18910_bits_payload_client_xact_id;
  assign gntNet_io_in_1_bits_payload_manager_xact_id = T_18910_bits_payload_manager_xact_id;
  assign gntNet_io_in_1_bits_payload_is_builtin_type = T_18910_bits_payload_is_builtin_type;
  assign gntNet_io_in_1_bits_payload_g_type = T_18910_bits_payload_g_type;
  assign gntNet_io_in_1_bits_payload_data = T_18910_bits_payload_data;
  assign gntNet_io_in_2_valid = 1'h0;
  assign gntNet_io_in_2_bits_header_src = GEN_42;
  assign gntNet_io_in_2_bits_header_dst = GEN_43;
  assign gntNet_io_in_2_bits_payload_addr_beat = GEN_44;
  assign gntNet_io_in_2_bits_payload_client_xact_id = GEN_45;
  assign gntNet_io_in_2_bits_payload_manager_xact_id = GEN_46;
  assign gntNet_io_in_2_bits_payload_is_builtin_type = GEN_47;
  assign gntNet_io_in_2_bits_payload_g_type = GEN_48;
  assign gntNet_io_in_2_bits_payload_data = GEN_49;
  assign gntNet_io_in_3_valid = 1'h0;
  assign gntNet_io_in_3_bits_header_src = GEN_50;
  assign gntNet_io_in_3_bits_header_dst = GEN_51;
  assign gntNet_io_in_3_bits_payload_addr_beat = GEN_52;
  assign gntNet_io_in_3_bits_payload_client_xact_id = GEN_53;
  assign gntNet_io_in_3_bits_payload_manager_xact_id = GEN_54;
  assign gntNet_io_in_3_bits_payload_is_builtin_type = GEN_55;
  assign gntNet_io_in_3_bits_payload_g_type = GEN_56;
  assign gntNet_io_in_3_bits_payload_data = GEN_57;
  assign gntNet_io_out_0_ready = 1'h0;
  assign gntNet_io_out_1_ready = 1'h0;
  assign gntNet_io_out_2_ready = T_19366_ready;
  assign gntNet_io_out_3_ready = T_20006_ready;
  assign ackNet_clk = clk;
  assign ackNet_reset = reset;
  assign ackNet_io_in_0_valid = 1'h0;
  assign ackNet_io_in_0_bits_header_src = GEN_58;
  assign ackNet_io_in_0_bits_header_dst = GEN_59;
  assign ackNet_io_in_0_bits_payload_manager_xact_id = GEN_60;
  assign ackNet_io_in_1_valid = 1'h0;
  assign ackNet_io_in_1_bits_header_src = GEN_61;
  assign ackNet_io_in_1_bits_header_dst = GEN_62;
  assign ackNet_io_in_1_bits_payload_manager_xact_id = GEN_63;
  assign ackNet_io_in_2_valid = T_21585_valid;
  assign ackNet_io_in_2_bits_header_src = T_21585_bits_header_src;
  assign ackNet_io_in_2_bits_header_dst = T_21585_bits_header_dst;
  assign ackNet_io_in_2_bits_payload_manager_xact_id = T_21585_bits_payload_manager_xact_id;
  assign ackNet_io_in_3_valid = T_21740_valid;
  assign ackNet_io_in_3_bits_header_src = T_21740_bits_header_src;
  assign ackNet_io_in_3_bits_header_dst = T_21740_bits_header_dst;
  assign ackNet_io_in_3_bits_payload_manager_xact_id = T_21740_bits_payload_manager_xact_id;
  assign ackNet_io_out_0_ready = T_20631_ready;
  assign ackNet_io_out_1_ready = T_21246_ready;
  assign ackNet_io_out_2_ready = 1'h0;
  assign ackNet_io_out_3_ready = 1'h0;
  assign T_14149_ready = TileLinkEnqueuer_2_1_io_client_acquire_ready;
  assign T_14149_valid = acqNet_io_out_0_valid;
  assign T_14149_bits_header_src = T_14408;
  assign T_14149_bits_header_dst = acqNet_io_out_0_bits_header_dst;
  assign T_14149_bits_payload_addr_block = acqNet_io_out_0_bits_payload_addr_block;
  assign T_14149_bits_payload_client_xact_id = acqNet_io_out_0_bits_payload_client_xact_id;
  assign T_14149_bits_payload_addr_beat = acqNet_io_out_0_bits_payload_addr_beat;
  assign T_14149_bits_payload_is_builtin_type = acqNet_io_out_0_bits_payload_is_builtin_type;
  assign T_14149_bits_payload_a_type = acqNet_io_out_0_bits_payload_a_type;
  assign T_14149_bits_payload_union = acqNet_io_out_0_bits_payload_union;
  assign T_14149_bits_payload_data = acqNet_io_out_0_bits_payload_data;
  assign T_14407 = acqNet_io_out_0_bits_header_src - 2'h2;
  assign T_14408 = T_14407[1:0];
  assign T_14794_ready = TileLinkEnqueuer_3_1_io_client_acquire_ready;
  assign T_14794_valid = acqNet_io_out_1_valid;
  assign T_14794_bits_header_src = T_15053;
  assign T_14794_bits_header_dst = acqNet_io_out_1_bits_header_dst;
  assign T_14794_bits_payload_addr_block = acqNet_io_out_1_bits_payload_addr_block;
  assign T_14794_bits_payload_client_xact_id = acqNet_io_out_1_bits_payload_client_xact_id;
  assign T_14794_bits_payload_addr_beat = acqNet_io_out_1_bits_payload_addr_beat;
  assign T_14794_bits_payload_is_builtin_type = acqNet_io_out_1_bits_payload_is_builtin_type;
  assign T_14794_bits_payload_a_type = acqNet_io_out_1_bits_payload_a_type;
  assign T_14794_bits_payload_union = acqNet_io_out_1_bits_payload_union;
  assign T_14794_bits_payload_data = acqNet_io_out_1_bits_payload_data;
  assign T_15052 = acqNet_io_out_1_bits_header_src - 2'h2;
  assign T_15053 = T_15052[1:0];
  assign T_15163_ready = acqNet_io_in_2_ready;
  assign T_15163_valid = TileLinkEnqueuer_4_io_manager_acquire_valid;
  assign T_15163_bits_header_src = T_15238;
  assign T_15163_bits_header_dst = TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  assign T_15163_bits_payload_addr_block = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  assign T_15163_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  assign T_15163_bits_payload_addr_beat = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  assign T_15163_bits_payload_is_builtin_type = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_15163_bits_payload_a_type = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  assign T_15163_bits_payload_union = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  assign T_15163_bits_payload_data = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  assign T_15237 = TileLinkEnqueuer_4_io_manager_acquire_bits_header_src + 2'h2;
  assign T_15238 = T_15237[1:0];
  assign T_15348_ready = acqNet_io_in_3_ready;
  assign T_15348_valid = TileLinkEnqueuer_1_1_io_manager_acquire_valid;
  assign T_15348_bits_header_src = T_15423;
  assign T_15348_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst;
  assign T_15348_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block;
  assign T_15348_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id;
  assign T_15348_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat;
  assign T_15348_bits_payload_is_builtin_type = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_15348_bits_payload_a_type = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type;
  assign T_15348_bits_payload_union = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union;
  assign T_15348_bits_payload_data = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data;
  assign T_15422 = TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src + 2'h2;
  assign T_15423 = T_15422[1:0];
  assign T_15806_ready = TileLinkEnqueuer_2_1_io_client_release_ready;
  assign T_15806_valid = relNet_io_out_0_valid;
  assign T_15806_bits_header_src = T_16063;
  assign T_15806_bits_header_dst = relNet_io_out_0_bits_header_dst;
  assign T_15806_bits_payload_addr_beat = relNet_io_out_0_bits_payload_addr_beat;
  assign T_15806_bits_payload_addr_block = relNet_io_out_0_bits_payload_addr_block;
  assign T_15806_bits_payload_client_xact_id = relNet_io_out_0_bits_payload_client_xact_id;
  assign T_15806_bits_payload_voluntary = relNet_io_out_0_bits_payload_voluntary;
  assign T_15806_bits_payload_r_type = relNet_io_out_0_bits_payload_r_type;
  assign T_15806_bits_payload_data = relNet_io_out_0_bits_payload_data;
  assign T_16062 = relNet_io_out_0_bits_header_src - 2'h2;
  assign T_16063 = T_16062[1:0];
  assign T_16446_ready = TileLinkEnqueuer_3_1_io_client_release_ready;
  assign T_16446_valid = relNet_io_out_1_valid;
  assign T_16446_bits_header_src = T_16703;
  assign T_16446_bits_header_dst = relNet_io_out_1_bits_header_dst;
  assign T_16446_bits_payload_addr_beat = relNet_io_out_1_bits_payload_addr_beat;
  assign T_16446_bits_payload_addr_block = relNet_io_out_1_bits_payload_addr_block;
  assign T_16446_bits_payload_client_xact_id = relNet_io_out_1_bits_payload_client_xact_id;
  assign T_16446_bits_payload_voluntary = relNet_io_out_1_bits_payload_voluntary;
  assign T_16446_bits_payload_r_type = relNet_io_out_1_bits_payload_r_type;
  assign T_16446_bits_payload_data = relNet_io_out_1_bits_payload_data;
  assign T_16702 = relNet_io_out_1_bits_header_src - 2'h2;
  assign T_16703 = T_16702[1:0];
  assign T_16810_ready = relNet_io_in_2_ready;
  assign T_16810_valid = TileLinkEnqueuer_4_io_manager_release_valid;
  assign T_16810_bits_header_src = T_16883;
  assign T_16810_bits_header_dst = TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  assign T_16810_bits_payload_addr_beat = TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  assign T_16810_bits_payload_addr_block = TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  assign T_16810_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  assign T_16810_bits_payload_voluntary = TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  assign T_16810_bits_payload_r_type = TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  assign T_16810_bits_payload_data = TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  assign T_16882 = TileLinkEnqueuer_4_io_manager_release_bits_header_src + 2'h2;
  assign T_16883 = T_16882[1:0];
  assign T_16990_ready = relNet_io_in_3_ready;
  assign T_16990_valid = TileLinkEnqueuer_1_1_io_manager_release_valid;
  assign T_16990_bits_header_src = T_17063;
  assign T_16990_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst;
  assign T_16990_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat;
  assign T_16990_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block;
  assign T_16990_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id;
  assign T_16990_bits_payload_voluntary = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary;
  assign T_16990_bits_payload_r_type = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type;
  assign T_16990_bits_payload_data = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data;
  assign T_17062 = TileLinkEnqueuer_1_1_io_manager_release_bits_header_src + 2'h2;
  assign T_17063 = T_17062[1:0];
  assign T_17158_ready = prbNet_io_in_0_ready;
  assign T_17158_valid = TileLinkEnqueuer_2_1_io_client_probe_valid;
  assign T_17158_bits_header_src = TileLinkEnqueuer_2_1_io_client_probe_bits_header_src;
  assign T_17158_bits_header_dst = T_17223;
  assign T_17158_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block;
  assign T_17158_bits_payload_p_type = TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type;
  assign T_17222 = TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst + 2'h2;
  assign T_17223 = T_17222[1:0];
  assign T_17318_ready = prbNet_io_in_1_ready;
  assign T_17318_valid = TileLinkEnqueuer_3_1_io_client_probe_valid;
  assign T_17318_bits_header_src = TileLinkEnqueuer_3_1_io_client_probe_bits_header_src;
  assign T_17318_bits_header_dst = T_17383;
  assign T_17318_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block;
  assign T_17318_bits_payload_p_type = TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type;
  assign T_17382 = TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst + 2'h2;
  assign T_17383 = T_17382[1:0];
  assign T_17754_ready = TileLinkEnqueuer_4_io_manager_probe_ready;
  assign T_17754_valid = prbNet_io_out_2_valid;
  assign T_17754_bits_header_src = prbNet_io_out_2_bits_header_src;
  assign T_17754_bits_header_dst = T_18003;
  assign T_17754_bits_payload_addr_block = prbNet_io_out_2_bits_payload_addr_block;
  assign T_17754_bits_payload_p_type = prbNet_io_out_2_bits_payload_p_type;
  assign T_18002 = prbNet_io_out_2_bits_header_dst - 2'h2;
  assign T_18003 = T_18002[1:0];
  assign T_18374_ready = TileLinkEnqueuer_1_1_io_manager_probe_ready;
  assign T_18374_valid = prbNet_io_out_3_valid;
  assign T_18374_bits_header_src = prbNet_io_out_3_bits_header_src;
  assign T_18374_bits_header_dst = T_18623;
  assign T_18374_bits_payload_addr_block = prbNet_io_out_3_bits_payload_addr_block;
  assign T_18374_bits_payload_p_type = prbNet_io_out_3_bits_payload_p_type;
  assign T_18622 = prbNet_io_out_3_bits_header_dst - 2'h2;
  assign T_18623 = T_18622[1:0];
  assign T_18730_ready = gntNet_io_in_0_ready;
  assign T_18730_valid = TileLinkEnqueuer_2_1_io_client_grant_valid;
  assign T_18730_bits_header_src = TileLinkEnqueuer_2_1_io_client_grant_bits_header_src;
  assign T_18730_bits_header_dst = T_18803;
  assign T_18730_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat;
  assign T_18730_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id;
  assign T_18730_bits_payload_manager_xact_id = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id;
  assign T_18730_bits_payload_is_builtin_type = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type;
  assign T_18730_bits_payload_g_type = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type;
  assign T_18730_bits_payload_data = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data;
  assign T_18802 = TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst + 2'h2;
  assign T_18803 = T_18802[1:0];
  assign T_18910_ready = gntNet_io_in_1_ready;
  assign T_18910_valid = TileLinkEnqueuer_3_1_io_client_grant_valid;
  assign T_18910_bits_header_src = TileLinkEnqueuer_3_1_io_client_grant_bits_header_src;
  assign T_18910_bits_header_dst = T_18983;
  assign T_18910_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat;
  assign T_18910_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id;
  assign T_18910_bits_payload_manager_xact_id = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id;
  assign T_18910_bits_payload_is_builtin_type = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type;
  assign T_18910_bits_payload_g_type = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type;
  assign T_18910_bits_payload_data = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data;
  assign T_18982 = TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst + 2'h2;
  assign T_18983 = T_18982[1:0];
  assign T_19366_ready = TileLinkEnqueuer_4_io_manager_grant_ready;
  assign T_19366_valid = gntNet_io_out_2_valid;
  assign T_19366_bits_header_src = gntNet_io_out_2_bits_header_src;
  assign T_19366_bits_header_dst = T_19623;
  assign T_19366_bits_payload_addr_beat = gntNet_io_out_2_bits_payload_addr_beat;
  assign T_19366_bits_payload_client_xact_id = gntNet_io_out_2_bits_payload_client_xact_id;
  assign T_19366_bits_payload_manager_xact_id = gntNet_io_out_2_bits_payload_manager_xact_id;
  assign T_19366_bits_payload_is_builtin_type = gntNet_io_out_2_bits_payload_is_builtin_type;
  assign T_19366_bits_payload_g_type = gntNet_io_out_2_bits_payload_g_type;
  assign T_19366_bits_payload_data = gntNet_io_out_2_bits_payload_data;
  assign T_19622 = gntNet_io_out_2_bits_header_dst - 2'h2;
  assign T_19623 = T_19622[1:0];
  assign T_20006_ready = TileLinkEnqueuer_1_1_io_manager_grant_ready;
  assign T_20006_valid = gntNet_io_out_3_valid;
  assign T_20006_bits_header_src = gntNet_io_out_3_bits_header_src;
  assign T_20006_bits_header_dst = T_20263;
  assign T_20006_bits_payload_addr_beat = gntNet_io_out_3_bits_payload_addr_beat;
  assign T_20006_bits_payload_client_xact_id = gntNet_io_out_3_bits_payload_client_xact_id;
  assign T_20006_bits_payload_manager_xact_id = gntNet_io_out_3_bits_payload_manager_xact_id;
  assign T_20006_bits_payload_is_builtin_type = gntNet_io_out_3_bits_payload_is_builtin_type;
  assign T_20006_bits_payload_g_type = gntNet_io_out_3_bits_payload_g_type;
  assign T_20006_bits_payload_data = gntNet_io_out_3_bits_payload_data;
  assign T_20262 = gntNet_io_out_3_bits_header_dst - 2'h2;
  assign T_20263 = T_20262[1:0];
  assign T_20631_ready = TileLinkEnqueuer_2_1_io_client_finish_ready;
  assign T_20631_valid = ackNet_io_out_0_valid;
  assign T_20631_bits_header_src = T_20878;
  assign T_20631_bits_header_dst = ackNet_io_out_0_bits_header_dst;
  assign T_20631_bits_payload_manager_xact_id = ackNet_io_out_0_bits_payload_manager_xact_id;
  assign T_20877 = ackNet_io_out_0_bits_header_src - 2'h2;
  assign T_20878 = T_20877[1:0];
  assign T_21246_ready = TileLinkEnqueuer_3_1_io_client_finish_ready;
  assign T_21246_valid = ackNet_io_out_1_valid;
  assign T_21246_bits_header_src = T_21493;
  assign T_21246_bits_header_dst = ackNet_io_out_1_bits_header_dst;
  assign T_21246_bits_payload_manager_xact_id = ackNet_io_out_1_bits_payload_manager_xact_id;
  assign T_21492 = ackNet_io_out_1_bits_header_src - 2'h2;
  assign T_21493 = T_21492[1:0];
  assign T_21585_ready = ackNet_io_in_2_ready;
  assign T_21585_valid = TileLinkEnqueuer_4_io_manager_finish_valid;
  assign T_21585_bits_header_src = T_21648;
  assign T_21585_bits_header_dst = TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  assign T_21585_bits_payload_manager_xact_id = TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  assign T_21647 = TileLinkEnqueuer_4_io_manager_finish_bits_header_src + 2'h2;
  assign T_21648 = T_21647[1:0];
  assign T_21740_ready = ackNet_io_in_3_ready;
  assign T_21740_valid = TileLinkEnqueuer_1_1_io_manager_finish_valid;
  assign T_21740_bits_header_src = T_21803;
  assign T_21740_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst;
  assign T_21740_bits_payload_manager_xact_id = TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id;
  assign T_21802 = TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src + 2'h2;
  assign T_21803 = T_21802[1:0];
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_64 = {1{$random}};
  GEN_0 = GEN_64[1:0];
  GEN_65 = {1{$random}};
  GEN_1 = GEN_65[1:0];
  GEN_66 = {1{$random}};
  GEN_2 = GEN_66[25:0];
  GEN_67 = {1{$random}};
  GEN_3 = GEN_67[1:0];
  GEN_68 = {1{$random}};
  GEN_4 = GEN_68[2:0];
  GEN_69 = {1{$random}};
  GEN_5 = GEN_69[0:0];
  GEN_70 = {1{$random}};
  GEN_6 = GEN_70[2:0];
  GEN_71 = {1{$random}};
  GEN_7 = GEN_71[11:0];
  GEN_72 = {2{$random}};
  GEN_8 = GEN_72[63:0];
  GEN_73 = {1{$random}};
  GEN_9 = GEN_73[1:0];
  GEN_74 = {1{$random}};
  GEN_10 = GEN_74[1:0];
  GEN_75 = {1{$random}};
  GEN_11 = GEN_75[25:0];
  GEN_76 = {1{$random}};
  GEN_12 = GEN_76[1:0];
  GEN_77 = {1{$random}};
  GEN_13 = GEN_77[2:0];
  GEN_78 = {1{$random}};
  GEN_14 = GEN_78[0:0];
  GEN_79 = {1{$random}};
  GEN_15 = GEN_79[2:0];
  GEN_80 = {1{$random}};
  GEN_16 = GEN_80[11:0];
  GEN_81 = {2{$random}};
  GEN_17 = GEN_81[63:0];
  GEN_82 = {1{$random}};
  GEN_18 = GEN_82[1:0];
  GEN_83 = {1{$random}};
  GEN_19 = GEN_83[1:0];
  GEN_84 = {1{$random}};
  GEN_20 = GEN_84[2:0];
  GEN_85 = {1{$random}};
  GEN_21 = GEN_85[25:0];
  GEN_86 = {1{$random}};
  GEN_22 = GEN_86[1:0];
  GEN_87 = {1{$random}};
  GEN_23 = GEN_87[0:0];
  GEN_88 = {1{$random}};
  GEN_24 = GEN_88[2:0];
  GEN_89 = {2{$random}};
  GEN_25 = GEN_89[63:0];
  GEN_90 = {1{$random}};
  GEN_26 = GEN_90[1:0];
  GEN_91 = {1{$random}};
  GEN_27 = GEN_91[1:0];
  GEN_92 = {1{$random}};
  GEN_28 = GEN_92[2:0];
  GEN_93 = {1{$random}};
  GEN_29 = GEN_93[25:0];
  GEN_94 = {1{$random}};
  GEN_30 = GEN_94[1:0];
  GEN_95 = {1{$random}};
  GEN_31 = GEN_95[0:0];
  GEN_96 = {1{$random}};
  GEN_32 = GEN_96[2:0];
  GEN_97 = {2{$random}};
  GEN_33 = GEN_97[63:0];
  GEN_98 = {1{$random}};
  GEN_34 = GEN_98[1:0];
  GEN_99 = {1{$random}};
  GEN_35 = GEN_99[1:0];
  GEN_100 = {1{$random}};
  GEN_36 = GEN_100[25:0];
  GEN_101 = {1{$random}};
  GEN_37 = GEN_101[1:0];
  GEN_102 = {1{$random}};
  GEN_38 = GEN_102[1:0];
  GEN_103 = {1{$random}};
  GEN_39 = GEN_103[1:0];
  GEN_104 = {1{$random}};
  GEN_40 = GEN_104[25:0];
  GEN_105 = {1{$random}};
  GEN_41 = GEN_105[1:0];
  GEN_106 = {1{$random}};
  GEN_42 = GEN_106[1:0];
  GEN_107 = {1{$random}};
  GEN_43 = GEN_107[1:0];
  GEN_108 = {1{$random}};
  GEN_44 = GEN_108[2:0];
  GEN_109 = {1{$random}};
  GEN_45 = GEN_109[1:0];
  GEN_110 = {1{$random}};
  GEN_46 = GEN_110[2:0];
  GEN_111 = {1{$random}};
  GEN_47 = GEN_111[0:0];
  GEN_112 = {1{$random}};
  GEN_48 = GEN_112[3:0];
  GEN_113 = {2{$random}};
  GEN_49 = GEN_113[63:0];
  GEN_114 = {1{$random}};
  GEN_50 = GEN_114[1:0];
  GEN_115 = {1{$random}};
  GEN_51 = GEN_115[1:0];
  GEN_116 = {1{$random}};
  GEN_52 = GEN_116[2:0];
  GEN_117 = {1{$random}};
  GEN_53 = GEN_117[1:0];
  GEN_118 = {1{$random}};
  GEN_54 = GEN_118[2:0];
  GEN_119 = {1{$random}};
  GEN_55 = GEN_119[0:0];
  GEN_120 = {1{$random}};
  GEN_56 = GEN_120[3:0];
  GEN_121 = {2{$random}};
  GEN_57 = GEN_121[63:0];
  GEN_122 = {1{$random}};
  GEN_58 = GEN_122[1:0];
  GEN_123 = {1{$random}};
  GEN_59 = GEN_123[1:0];
  GEN_124 = {1{$random}};
  GEN_60 = GEN_124[2:0];
  GEN_125 = {1{$random}};
  GEN_61 = GEN_125[1:0];
  GEN_126 = {1{$random}};
  GEN_62 = GEN_126[1:0];
  GEN_127 = {1{$random}};
  GEN_63 = GEN_127[2:0];
  end
`endif
endmodule
module BufferedBroadcastVoluntaryReleaseTracker(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should
);
  wire  T_44;
  reg [3:0] T_55;
  reg [31:0] GEN_28;
  reg [25:0] T_57;
  reg [31:0] GEN_29;
  reg [2:0] T_59;
  reg [31:0] GEN_30;
  reg  T_61;
  reg [31:0] GEN_31;
  reg [1:0] T_63;
  reg [31:0] GEN_32;
  reg [7:0] T_65;
  reg [31:0] GEN_33;
  wire  T_74_pending;
  wire [2:0] T_74_up_idx;
  wire  T_74_up_done;
  wire [2:0] T_74_down_idx;
  wire  T_74_down_done;
  reg  T_83;
  reg [31:0] GEN_35;
  reg [7:0] T_85;
  reg [31:0] GEN_36;
  wire  T_94_pending;
  wire [2:0] T_94_up_idx;
  wire  T_94_up_done;
  wire [2:0] T_94_down_idx;
  wire  T_94_down_done;
  wire [7:0] GEN_76;
  wire  T_103;
  wire  T_104;
  wire  T_105;
  wire  T_131_sharers;
  wire [1:0] T_183_state;
  wire  T_279_inner_sharers;
  wire [1:0] T_279_outer_state;
  wire  T_1617;
  wire  T_1618;
  wire  T_1619;
  wire  T_1620;
  wire  T_1622;
  wire  T_1623;
  wire  T_1625;
  wire  T_1626;
  wire  T_1628;
  wire [63:0] T_1642_0;
  wire [63:0] T_1642_1;
  wire [63:0] T_1642_2;
  wire [63:0] T_1642_3;
  wire [63:0] T_1642_4;
  wire [63:0] T_1642_5;
  wire [63:0] T_1642_6;
  wire [63:0] T_1642_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_37;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_46;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_55;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_56;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_57;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_58;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_59;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_60;
  wire  T_1647;
  wire  T_1648;
  wire  T_1649;
  wire  T_1651;
  wire  T_1652;
  wire  T_1654;
  wire  T_1655;
  wire  T_1660;
  wire  T_1664;
  wire  T_1665;
  wire  T_1670;
  wire [2:0] T_1677_0;
  wire [2:0] T_1677_1;
  wire [2:0] T_1677_2;
  wire  T_1679;
  wire  T_1680;
  wire  T_1681;
  wire  T_1684;
  wire  T_1685;
  wire  T_1687;
  reg [2:0] T_1689;
  reg [31:0] GEN_82;
  wire  T_1691;
  wire [2:0] GEN_77;
  wire [3:0] T_1693;
  wire [2:0] T_1694;
  wire [2:0] GEN_2;
  wire  T_1695;
  wire [2:0] T_1696;
  wire  T_1697;
  wire  T_1698;
  wire [3:0] GEN_78;
  wire  T_1701;
  wire  T_1702;
  wire  T_1703;
  wire  T_1704;
  wire [2:0] T_1712_0;
  wire [3:0] GEN_79;
  wire  T_1714;
  wire [1:0] T_1722_0;
  wire [1:0] T_1722_1;
  wire [3:0] GEN_80;
  wire  T_1724;
  wire [3:0] GEN_81;
  wire  T_1725;
  wire  T_1728;
  wire  T_1729;
  wire  T_1731;
  reg [2:0] T_1733;
  reg [31:0] GEN_86;
  wire  T_1735;
  wire [3:0] T_1737;
  wire [2:0] T_1738;
  wire [2:0] GEN_3;
  wire  T_1739;
  wire [2:0] T_1740;
  wire  T_1741;
  reg  T_1743;
  reg [31:0] GEN_88;
  wire  T_1745;
  wire  T_1746;
  wire [1:0] T_1748;
  wire  T_1749;
  wire  GEN_4;
  wire  T_1751;
  wire  T_1752;
  wire [1:0] T_1754;
  wire  T_1755;
  wire  GEN_5;
  wire  T_1757;
  wire  T_1759;
  wire  T_1760;
  wire [25:0] GEN_6;
  wire [3:0] GEN_7;
  wire [2:0] T_1769_0;
  wire [2:0] T_1769_1;
  wire [2:0] T_1769_2;
  wire [2:0] GEN_83;
  wire [2:0] T_1792_0;
  wire [2:0] T_1792_1;
  wire [2:0] T_1792_2;
  wire  T_1794;
  wire  T_1795;
  wire  T_1796;
  wire  T_1799;
  wire  T_1800;
  wire [2:0] T_1808_0;
  wire [2:0] T_1808_1;
  wire [2:0] T_1808_2;
  wire  T_1810;
  wire  T_1811;
  wire  T_1812;
  wire  T_1815;
  wire  T_1816;
  wire  T_1817;
  wire [7:0] GEN_84;
  wire [8:0] T_1819;
  wire [7:0] T_1820;
  wire [7:0] T_1821;
  wire [7:0] GEN_85;
  wire [7:0] T_1823;
  wire [7:0] T_1824;
  wire [7:0] T_1825;
  wire [7:0] T_1827;
  wire [2:0] GEN_8;
  wire  GEN_9;
  wire [1:0] GEN_10;
  wire [7:0] GEN_17;
  wire  T_1829;
  wire  T_1831;
  wire  T_1832;
  wire  T_1834;
  wire  T_1835;
  wire [2:0] T_1842_0;
  wire [2:0] T_1842_1;
  wire [2:0] T_1842_2;
  wire  T_1844;
  wire  T_1845;
  wire  T_1846;
  wire  T_1849;
  wire  T_1850;
  wire  T_1851;
  wire [7:0] GEN_87;
  wire [8:0] T_1853;
  wire [7:0] T_1854;
  wire [7:0] T_1855;
  wire [7:0] T_1859;
  wire [7:0] T_1860;
  wire [7:0] GEN_21;
  wire [2:0] GEN_25;
  wire  GEN_26;
  wire [1:0] GEN_27;
  wire [7:0] GEN_34;
  wire [3:0] T_1866_0;
  wire [3:0] T_1866_1;
  wire [3:0] T_1866_2;
  wire [3:0] T_1866_3;
  wire  T_1868;
  wire  T_1869;
  wire  T_1870;
  wire  T_1871;
  wire  T_1874;
  wire  T_1875;
  wire  T_1876;
  wire  T_1877;
  wire  T_1880;
  wire  T_1882;
  wire  T_1883;
  wire [2:0] T_1918_addr_beat;
  wire [25:0] T_1918_addr_block;
  wire [1:0] T_1918_client_xact_id;
  wire  T_1918_voluntary;
  wire [2:0] T_1918_r_type;
  wire [63:0] T_1918_data;
  wire  T_1918_client_id;
  wire [2:0] T_1985_addr_beat;
  wire [1:0] T_1985_client_xact_id;
  wire [2:0] T_1985_manager_xact_id;
  wire  T_1985_is_builtin_type;
  wire [3:0] T_1985_g_type;
  wire [63:0] T_1985_data;
  wire  T_1985_client_id;
  wire  T_2026;
  wire [63:0] GEN_0;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  wire [2:0] GEN_94;
  wire [63:0] GEN_40;
  wire [2:0] GEN_95;
  wire [63:0] GEN_41;
  wire [63:0] GEN_42;
  wire [63:0] GEN_43;
  wire [63:0] GEN_44;
  wire [63:0] GEN_45;
  wire [63:0] GEN_47;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  wire [63:0] GEN_50;
  wire [63:0] GEN_51;
  wire [63:0] GEN_52;
  wire [63:0] GEN_53;
  wire [63:0] GEN_54;
  wire [1:0] T_2058_state;
  wire  T_2086;
  wire  T_2087;
  wire [2:0] T_2093_0;
  wire [2:0] T_2093_1;
  wire [2:0] T_2093_2;
  wire  T_2095;
  wire  T_2096;
  wire  T_2097;
  wire  T_2100;
  wire  T_2101;
  wire  T_2102;
  wire [7:0] GEN_96;
  wire [8:0] T_2104;
  wire [7:0] T_2105;
  wire [7:0] T_2106;
  wire [7:0] T_2108;
  wire [7:0] T_2109;
  wire [7:0] T_2110;
  wire [7:0] T_2111;
  wire [2:0] T_2119_0;
  wire [2:0] T_2119_1;
  wire [2:0] T_2119_2;
  wire  T_2121;
  wire  T_2122;
  wire  T_2123;
  wire  T_2126;
  wire  T_2127;
  wire  T_2128;
  wire [7:0] GEN_98;
  wire [8:0] T_2131;
  wire [7:0] T_2132;
  wire [7:0] T_2135;
  wire [7:0] T_2136;
  wire [7:0] T_2137;
  wire [7:0] GEN_61;
  wire  GEN_62;
  wire  GEN_63;
  wire  T_2147;
  wire [2:0] T_2154_0;
  wire [2:0] T_2154_1;
  wire [2:0] T_2154_2;
  wire  T_2156;
  wire  T_2157;
  wire  T_2158;
  wire  T_2161;
  wire  T_2162;
  wire  T_2164;
  reg [2:0] T_2166;
  reg [31:0] GEN_89;
  wire  T_2168;
  wire [3:0] T_2170;
  wire [2:0] T_2171;
  wire [2:0] GEN_64;
  wire  T_2172;
  wire [2:0] T_2173;
  wire  T_2174;
  wire  T_2175;
  wire  T_2177;
  wire  T_2178;
  wire  T_2179;
  wire [2:0] T_2187_0;
  wire [3:0] GEN_103;
  wire  T_2189;
  wire  T_2197_0;
  wire [3:0] GEN_104;
  wire  T_2199;
  wire  T_2202;
  wire  T_2204;
  reg [2:0] T_2206;
  reg [31:0] GEN_90;
  wire  T_2208;
  wire [3:0] T_2210;
  wire [2:0] T_2211;
  wire [2:0] GEN_65;
  wire  T_2212;
  wire [2:0] T_2213;
  wire  T_2214;
  reg  T_2216;
  reg [31:0] GEN_91;
  wire  T_2218;
  wire  T_2219;
  wire [1:0] T_2221;
  wire  T_2222;
  wire  GEN_66;
  wire  T_2224;
  wire  T_2225;
  wire [1:0] T_2227;
  wire  T_2228;
  wire  GEN_67;
  wire  T_2230;
  wire  T_2231;
  wire [2:0] T_2237_0;
  wire [2:0] T_2237_1;
  wire [2:0] T_2237_2;
  wire  T_2239;
  wire  T_2240;
  wire  T_2241;
  wire  T_2244;
  wire  T_2245;
  wire [7:0] T_2246;
  wire  T_2247;
  wire  T_2249;
  wire  T_2250;
  wire [1:0] T_2258_0;
  wire  T_2260;
  wire [2:0] T_2263;
  wire [2:0] T_2299_addr_beat;
  wire [25:0] T_2299_addr_block;
  wire [2:0] T_2299_client_xact_id;
  wire  T_2299_voluntary;
  wire [2:0] T_2299_r_type;
  wire [63:0] T_2299_data;
  wire [63:0] GEN_1;
  wire [63:0] GEN_68;
  wire [63:0] GEN_69;
  wire [63:0] GEN_70;
  wire [63:0] GEN_71;
  wire [63:0] GEN_72;
  wire [63:0] GEN_73;
  wire [63:0] GEN_74;
  wire  T_2329;
  wire  T_2330;
  wire  T_2331;
  wire  T_2333;
  wire  T_2335;
  wire [3:0] GEN_75;
  reg [25:0] GEN_11;
  reg [31:0] GEN_92;
  reg [1:0] GEN_12;
  reg [31:0] GEN_93;
  reg  GEN_13;
  reg [31:0] GEN_97;
  reg [25:0] GEN_14;
  reg [31:0] GEN_99;
  reg [2:0] GEN_15;
  reg [31:0] GEN_100;
  reg [2:0] GEN_16;
  reg [31:0] GEN_101;
  reg  GEN_18;
  reg [31:0] GEN_102;
  reg [2:0] GEN_19;
  reg [31:0] GEN_105;
  reg [11:0] GEN_20;
  reg [31:0] GEN_106;
  reg [63:0] GEN_22;
  reg [63:0] GEN_107;
  reg  GEN_23;
  reg [31:0] GEN_108;
  reg  GEN_24;
  reg [31:0] GEN_109;
  assign io_inner_acquire_ready = 1'h0;
  assign io_inner_grant_valid = T_1883;
  assign io_inner_grant_bits_addr_beat = T_1985_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_1985_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = T_1985_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = T_1985_is_builtin_type;
  assign io_inner_grant_bits_g_type = T_1985_g_type;
  assign io_inner_grant_bits_data = T_1985_data;
  assign io_inner_grant_bits_client_id = T_1985_client_id;
  assign io_inner_finish_ready = 1'h0;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_11;
  assign io_inner_probe_bits_p_type = GEN_12;
  assign io_inner_probe_bits_client_id = GEN_13;
  assign io_inner_release_ready = T_2026;
  assign io_outer_acquire_valid = 1'h0;
  assign io_outer_acquire_bits_addr_block = GEN_14;
  assign io_outer_acquire_bits_client_xact_id = GEN_15;
  assign io_outer_acquire_bits_addr_beat = GEN_16;
  assign io_outer_acquire_bits_is_builtin_type = GEN_18;
  assign io_outer_acquire_bits_a_type = GEN_19;
  assign io_outer_acquire_bits_union = GEN_20;
  assign io_outer_acquire_bits_data = GEN_22;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2250;
  assign io_outer_release_bits_addr_beat = T_2299_addr_beat;
  assign io_outer_release_bits_addr_block = T_2299_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2299_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2299_voluntary;
  assign io_outer_release_bits_r_type = T_2299_r_type;
  assign io_outer_release_bits_data = T_2299_data;
  assign io_outer_grant_ready = T_2231;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_23;
  assign io_outer_finish_bits_manager_id = GEN_24;
  assign io_alloc_iacq_matches = T_1649;
  assign io_alloc_iacq_can = 1'h0;
  assign io_alloc_irel_matches = T_1652;
  assign io_alloc_irel_can = T_1617;
  assign io_alloc_oprb_matches = T_1655;
  assign io_alloc_oprb_can = 1'h0;
  assign T_44 = T_2333;
  assign T_74_pending = T_1757;
  assign T_74_up_idx = T_1696;
  assign T_74_up_done = T_1697;
  assign T_74_down_idx = T_1740;
  assign T_74_down_done = T_1741;
  assign T_94_pending = T_2230;
  assign T_94_up_idx = T_2173;
  assign T_94_up_done = T_2174;
  assign T_94_down_idx = T_2213;
  assign T_94_down_done = T_2214;
  assign GEN_76 = {{7'd0}, 1'h0};
  assign T_103 = T_85 != GEN_76;
  assign T_104 = T_83 | T_103;
  assign T_105 = T_104 | T_94_pending;
  assign T_131_sharers = 1'h0;
  assign T_183_state = {{1'd0}, 1'h0};
  assign T_279_inner_sharers = T_131_sharers;
  assign T_279_outer_state = T_183_state;
  assign T_1617 = T_55 == 4'h0;
  assign T_1618 = io_inner_release_ready & io_inner_release_valid;
  assign T_1619 = T_1617 & T_1618;
  assign T_1620 = T_1619 & io_alloc_irel_should;
  assign T_1622 = io_inner_release_bits_voluntary == 1'h0;
  assign T_1623 = T_1620 & T_1622;
  assign T_1625 = T_1623 == 1'h0;
  assign T_1626 = T_1625 | reset;
  assign T_1628 = T_1626 == 1'h0;
  assign T_1642_0 = 64'h0;
  assign T_1642_1 = 64'h0;
  assign T_1642_2 = 64'h0;
  assign T_1642_3 = 64'h0;
  assign T_1642_4 = 64'h0;
  assign T_1642_5 = 64'h0;
  assign T_1642_6 = 64'h0;
  assign T_1642_7 = 64'h0;
  assign T_1647 = T_55 != 4'h0;
  assign T_1648 = io_inner_acquire_bits_addr_block == T_57;
  assign T_1649 = T_1647 & T_1648;
  assign T_1651 = io_inner_release_bits_addr_block == T_57;
  assign T_1652 = T_1647 & T_1651;
  assign T_1654 = io_outer_probe_bits_addr_block == T_57;
  assign T_1655 = T_1647 & T_1654;
  assign T_1660 = T_105 | T_94_pending;
  assign T_1664 = T_1617 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_1665 = T_1664 & io_inner_release_bits_voluntary;
  assign T_1670 = T_1618 & T_1665;
  assign T_1677_0 = 3'h0;
  assign T_1677_1 = 3'h1;
  assign T_1677_2 = 3'h2;
  assign T_1679 = T_1677_0 == io_inner_release_bits_r_type;
  assign T_1680 = T_1677_1 == io_inner_release_bits_r_type;
  assign T_1681 = T_1677_2 == io_inner_release_bits_r_type;
  assign T_1684 = T_1679 | T_1680;
  assign T_1685 = T_1684 | T_1681;
  assign T_1687 = T_1670 & T_1685;
  assign T_1691 = T_1689 == 3'h7;
  assign GEN_77 = {{2'd0}, 1'h1};
  assign T_1693 = T_1689 + GEN_77;
  assign T_1694 = T_1693[2:0];
  assign GEN_2 = T_1687 ? T_1694 : T_1689;
  assign T_1695 = T_1687 & T_1691;
  assign T_1696 = T_1685 ? T_1689 : {{2'd0}, 1'h0};
  assign T_1697 = T_1685 ? T_1695 : T_1670;
  assign T_1698 = io_inner_grant_ready & io_inner_grant_valid;
  assign GEN_78 = {{1'd0}, 3'h0};
  assign T_1701 = io_inner_grant_bits_g_type == GEN_78;
  assign T_1702 = io_inner_grant_bits_is_builtin_type & T_1701;
  assign T_1703 = T_1647 & T_1702;
  assign T_1704 = T_1698 & T_1703;
  assign T_1712_0 = 3'h5;
  assign GEN_79 = {{1'd0}, T_1712_0};
  assign T_1714 = GEN_79 == io_inner_grant_bits_g_type;
  assign T_1722_0 = 2'h0;
  assign T_1722_1 = 2'h1;
  assign GEN_80 = {{2'd0}, T_1722_0};
  assign T_1724 = GEN_80 == io_inner_grant_bits_g_type;
  assign GEN_81 = {{2'd0}, T_1722_1};
  assign T_1725 = GEN_81 == io_inner_grant_bits_g_type;
  assign T_1728 = T_1724 | T_1725;
  assign T_1729 = io_inner_grant_bits_is_builtin_type ? T_1714 : T_1728;
  assign T_1731 = T_1704 & T_1729;
  assign T_1735 = T_1733 == 3'h7;
  assign T_1737 = T_1733 + GEN_77;
  assign T_1738 = T_1737[2:0];
  assign GEN_3 = T_1731 ? T_1738 : T_1733;
  assign T_1739 = T_1731 & T_1735;
  assign T_1740 = T_1729 ? T_1733 : {{2'd0}, 1'h0};
  assign T_1741 = T_1729 ? T_1739 : T_1704;
  assign T_1745 = T_1741 == 1'h0;
  assign T_1746 = T_1697 & T_1745;
  assign T_1748 = T_1743 + 1'h1;
  assign T_1749 = T_1748[0:0];
  assign GEN_4 = T_1746 ? T_1749 : T_1743;
  assign T_1751 = T_1697 == 1'h0;
  assign T_1752 = T_1741 & T_1751;
  assign T_1754 = T_1743 - 1'h1;
  assign T_1755 = T_1754[0:0];
  assign GEN_5 = T_1752 ? T_1755 : GEN_4;
  assign T_1757 = T_1743 > 1'h0;
  assign T_1759 = T_1617 & io_alloc_irel_should;
  assign T_1760 = T_1759 & io_inner_release_valid;
  assign GEN_6 = T_1760 ? io_inner_release_bits_addr_block : T_57;
  assign GEN_7 = T_1760 ? 4'h7 : T_55;
  assign T_1769_0 = 3'h0;
  assign T_1769_1 = 3'h1;
  assign T_1769_2 = 3'h2;
  assign GEN_83 = {{2'd0}, 1'h0};
  assign T_1792_0 = 3'h0;
  assign T_1792_1 = 3'h1;
  assign T_1792_2 = 3'h2;
  assign T_1794 = T_1792_0 == io_inner_release_bits_r_type;
  assign T_1795 = T_1792_1 == io_inner_release_bits_r_type;
  assign T_1796 = T_1792_2 == io_inner_release_bits_r_type;
  assign T_1799 = T_1794 | T_1795;
  assign T_1800 = T_1799 | T_1796;
  assign T_1808_0 = 3'h0;
  assign T_1808_1 = 3'h1;
  assign T_1808_2 = 3'h2;
  assign T_1810 = T_1808_0 == io_inner_release_bits_r_type;
  assign T_1811 = T_1808_1 == io_inner_release_bits_r_type;
  assign T_1812 = T_1808_2 == io_inner_release_bits_r_type;
  assign T_1815 = T_1810 | T_1811;
  assign T_1816 = T_1815 | T_1812;
  assign T_1817 = T_1618 & T_1816;
  assign GEN_84 = {{7'd0}, T_1817};
  assign T_1819 = 8'h0 - GEN_84;
  assign T_1820 = T_1819[7:0];
  assign T_1821 = ~ T_1820;
  assign GEN_85 = {{7'd0}, 1'h1};
  assign T_1823 = GEN_85 << io_inner_release_bits_addr_beat;
  assign T_1824 = ~ T_1823;
  assign T_1825 = T_1821 | T_1824;
  assign T_1827 = T_1800 ? T_1825 : {{7'd0}, 1'h0};
  assign GEN_8 = io_alloc_irel_should ? io_inner_release_bits_r_type : T_59;
  assign GEN_9 = io_alloc_irel_should ? io_inner_release_bits_client_id : T_61;
  assign GEN_10 = io_alloc_irel_should ? io_inner_release_bits_client_xact_id : T_63;
  assign GEN_17 = io_alloc_irel_should ? T_1827 : T_65;
  assign T_1829 = T_1651 & io_inner_release_bits_voluntary;
  assign T_1831 = T_65 != GEN_76;
  assign T_1832 = T_1829 & T_1831;
  assign T_1834 = io_alloc_irel_should == 1'h0;
  assign T_1835 = T_1834 & T_1832;
  assign T_1842_0 = 3'h0;
  assign T_1842_1 = 3'h1;
  assign T_1842_2 = 3'h2;
  assign T_1844 = T_1842_0 == io_inner_release_bits_r_type;
  assign T_1845 = T_1842_1 == io_inner_release_bits_r_type;
  assign T_1846 = T_1842_2 == io_inner_release_bits_r_type;
  assign T_1849 = T_1844 | T_1845;
  assign T_1850 = T_1849 | T_1846;
  assign T_1851 = T_1618 & T_1850;
  assign GEN_87 = {{7'd0}, T_1851};
  assign T_1853 = 8'h0 - GEN_87;
  assign T_1854 = T_1853[7:0];
  assign T_1855 = ~ T_1854;
  assign T_1859 = T_1855 | T_1824;
  assign T_1860 = T_65 & T_1859;
  assign GEN_21 = T_1835 ? T_1860 : GEN_17;
  assign GEN_25 = T_1618 ? GEN_8 : T_59;
  assign GEN_26 = T_1618 ? GEN_9 : T_61;
  assign GEN_27 = T_1618 ? GEN_10 : T_63;
  assign GEN_34 = T_1618 ? GEN_21 : T_65;
  assign T_1866_0 = 4'h3;
  assign T_1866_1 = 4'h4;
  assign T_1866_2 = 4'h5;
  assign T_1866_3 = 4'h7;
  assign T_1868 = T_1866_0 == T_55;
  assign T_1869 = T_1866_1 == T_55;
  assign T_1870 = T_1866_2 == T_55;
  assign T_1871 = T_1866_3 == T_55;
  assign T_1874 = T_1868 | T_1869;
  assign T_1875 = T_1874 | T_1870;
  assign T_1876 = T_1875 | T_1871;
  assign T_1877 = T_1876 & T_74_pending;
  assign T_1880 = T_1831 | T_1660;
  assign T_1882 = T_1880 == 1'h0;
  assign T_1883 = T_1877 & T_1882;
  assign T_1918_addr_beat = {{2'd0}, 1'h0};
  assign T_1918_addr_block = T_57;
  assign T_1918_client_xact_id = T_63;
  assign T_1918_voluntary = 1'h1;
  assign T_1918_r_type = T_59;
  assign T_1918_data = {{63'd0}, 1'h0};
  assign T_1918_client_id = T_61;
  assign T_1985_addr_beat = {{2'd0}, 1'h0};
  assign T_1985_client_xact_id = T_1918_client_xact_id;
  assign T_1985_manager_xact_id = {{2'd0}, 1'h0};
  assign T_1985_is_builtin_type = 1'h1;
  assign T_1985_g_type = {{1'd0}, 3'h0};
  assign T_1985_data = {{63'd0}, 1'h0};
  assign T_1985_client_id = T_1918_client_id;
  assign T_2026 = T_1617 | T_1832;
  assign GEN_0 = io_inner_release_bits_data;
  assign GEN_38 = GEN_83 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_0;
  assign GEN_39 = GEN_77 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_1;
  assign GEN_94 = {{1'd0}, 2'h2};
  assign GEN_40 = GEN_94 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_2;
  assign GEN_95 = {{1'd0}, 2'h3};
  assign GEN_41 = GEN_95 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_3;
  assign GEN_42 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_4;
  assign GEN_43 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_5;
  assign GEN_44 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_6;
  assign GEN_45 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_7;
  assign GEN_47 = T_1618 ? GEN_38 : data_buffer_0;
  assign GEN_48 = T_1618 ? GEN_39 : data_buffer_1;
  assign GEN_49 = T_1618 ? GEN_40 : data_buffer_2;
  assign GEN_50 = T_1618 ? GEN_41 : data_buffer_3;
  assign GEN_51 = T_1618 ? GEN_42 : data_buffer_4;
  assign GEN_52 = T_1618 ? GEN_43 : data_buffer_5;
  assign GEN_53 = T_1618 ? GEN_44 : data_buffer_6;
  assign GEN_54 = T_1618 ? GEN_45 : data_buffer_7;
  assign T_2058_state = 2'h2;
  assign T_2086 = T_1647 | io_alloc_irel_should;
  assign T_2087 = io_outer_release_ready & io_outer_release_valid;
  assign T_2093_0 = 3'h0;
  assign T_2093_1 = 3'h1;
  assign T_2093_2 = 3'h2;
  assign T_2095 = T_2093_0 == io_outer_release_bits_r_type;
  assign T_2096 = T_2093_1 == io_outer_release_bits_r_type;
  assign T_2097 = T_2093_2 == io_outer_release_bits_r_type;
  assign T_2100 = T_2095 | T_2096;
  assign T_2101 = T_2100 | T_2097;
  assign T_2102 = T_2087 & T_2101;
  assign GEN_96 = {{7'd0}, T_2102};
  assign T_2104 = 8'h0 - GEN_96;
  assign T_2105 = T_2104[7:0];
  assign T_2106 = ~ T_2105;
  assign T_2108 = GEN_85 << io_outer_release_bits_addr_beat;
  assign T_2109 = ~ T_2108;
  assign T_2110 = T_2106 | T_2109;
  assign T_2111 = T_85 & T_2110;
  assign T_2119_0 = 3'h0;
  assign T_2119_1 = 3'h1;
  assign T_2119_2 = 3'h2;
  assign T_2121 = T_2119_0 == io_inner_release_bits_r_type;
  assign T_2122 = T_2119_1 == io_inner_release_bits_r_type;
  assign T_2123 = T_2119_2 == io_inner_release_bits_r_type;
  assign T_2126 = T_2121 | T_2122;
  assign T_2127 = T_2126 | T_2123;
  assign T_2128 = T_1618 & T_2127;
  assign GEN_98 = {{7'd0}, T_2128};
  assign T_2131 = 8'h0 - GEN_98;
  assign T_2132 = T_2131[7:0];
  assign T_2135 = T_2132 & T_1823;
  assign T_2136 = T_2111 | T_2135;
  assign T_2137 = T_2136 | GEN_76;
  assign GEN_61 = T_2086 ? T_2137 : T_85;
  assign GEN_62 = T_1760 ? 1'h1 : T_83;
  assign GEN_63 = T_2087 ? 1'h0 : GEN_62;
  assign T_2147 = T_2087 & io_outer_release_bits_voluntary;
  assign T_2154_0 = 3'h0;
  assign T_2154_1 = 3'h1;
  assign T_2154_2 = 3'h2;
  assign T_2156 = T_2154_0 == io_outer_release_bits_r_type;
  assign T_2157 = T_2154_1 == io_outer_release_bits_r_type;
  assign T_2158 = T_2154_2 == io_outer_release_bits_r_type;
  assign T_2161 = T_2156 | T_2157;
  assign T_2162 = T_2161 | T_2158;
  assign T_2164 = T_2147 & T_2162;
  assign T_2168 = T_2166 == 3'h7;
  assign T_2170 = T_2166 + GEN_77;
  assign T_2171 = T_2170[2:0];
  assign GEN_64 = T_2164 ? T_2171 : T_2166;
  assign T_2172 = T_2164 & T_2168;
  assign T_2173 = T_2162 ? T_2166 : {{2'd0}, 1'h0};
  assign T_2174 = T_2162 ? T_2172 : T_2147;
  assign T_2175 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2177 = io_outer_grant_bits_g_type == GEN_78;
  assign T_2178 = io_outer_grant_bits_is_builtin_type & T_2177;
  assign T_2179 = T_2175 & T_2178;
  assign T_2187_0 = 3'h5;
  assign GEN_103 = {{1'd0}, T_2187_0};
  assign T_2189 = GEN_103 == io_outer_grant_bits_g_type;
  assign T_2197_0 = 1'h0;
  assign GEN_104 = {{3'd0}, T_2197_0};
  assign T_2199 = GEN_104 == io_outer_grant_bits_g_type;
  assign T_2202 = io_outer_grant_bits_is_builtin_type ? T_2189 : T_2199;
  assign T_2204 = T_2179 & T_2202;
  assign T_2208 = T_2206 == 3'h7;
  assign T_2210 = T_2206 + GEN_77;
  assign T_2211 = T_2210[2:0];
  assign GEN_65 = T_2204 ? T_2211 : T_2206;
  assign T_2212 = T_2204 & T_2208;
  assign T_2213 = T_2202 ? T_2206 : {{2'd0}, 1'h0};
  assign T_2214 = T_2202 ? T_2212 : T_2179;
  assign T_2218 = T_2214 == 1'h0;
  assign T_2219 = T_2174 & T_2218;
  assign T_2221 = T_2216 + 1'h1;
  assign T_2222 = T_2221[0:0];
  assign GEN_66 = T_2219 ? T_2222 : T_2216;
  assign T_2224 = T_2174 == 1'h0;
  assign T_2225 = T_2214 & T_2224;
  assign T_2227 = T_2216 - 1'h1;
  assign T_2228 = T_2227[0:0];
  assign GEN_67 = T_2225 ? T_2228 : GEN_66;
  assign T_2230 = T_2216 > 1'h0;
  assign T_2231 = T_55 == 4'h7;
  assign T_2237_0 = 3'h0;
  assign T_2237_1 = 3'h1;
  assign T_2237_2 = 3'h2;
  assign T_2239 = T_2237_0 == io_outer_release_bits_r_type;
  assign T_2240 = T_2237_1 == io_outer_release_bits_r_type;
  assign T_2241 = T_2237_2 == io_outer_release_bits_r_type;
  assign T_2244 = T_2239 | T_2240;
  assign T_2245 = T_2244 | T_2241;
  assign T_2246 = T_85 >> T_94_up_idx;
  assign T_2247 = T_2246[0];
  assign T_2249 = T_2245 ? T_2247 : T_105;
  assign T_2250 = T_2231 & T_2249;
  assign T_2258_0 = 2'h2;
  assign T_2260 = T_2258_0 == T_2058_state;
  assign T_2263 = T_2260 ? 3'h0 : 3'h3;
  assign T_2299_addr_beat = T_94_up_idx;
  assign T_2299_addr_block = T_57;
  assign T_2299_client_xact_id = {{2'd0}, 1'h0};
  assign T_2299_voluntary = 1'h1;
  assign T_2299_r_type = T_2263;
  assign T_2299_data = GEN_1;
  assign GEN_1 = GEN_74;
  assign GEN_68 = GEN_77 == T_94_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_69 = GEN_94 == T_94_up_idx ? data_buffer_2 : GEN_68;
  assign GEN_70 = GEN_95 == T_94_up_idx ? data_buffer_3 : GEN_69;
  assign GEN_71 = 3'h4 == T_94_up_idx ? data_buffer_4 : GEN_70;
  assign GEN_72 = 3'h5 == T_94_up_idx ? data_buffer_5 : GEN_71;
  assign GEN_73 = 3'h6 == T_94_up_idx ? data_buffer_6 : GEN_72;
  assign GEN_74 = 3'h7 == T_94_up_idx ? data_buffer_7 : GEN_73;
  assign T_2329 = T_1831 | T_74_pending;
  assign T_2330 = T_2329 | T_105;
  assign T_2331 = T_2330 | T_94_pending;
  assign T_2333 = T_2331 == 1'h0;
  assign T_2335 = T_2231 & T_44;
  assign GEN_75 = T_2335 ? 4'h0 : GEN_7;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_28 = {1{$random}};
  T_55 = GEN_28[3:0];
  GEN_29 = {1{$random}};
  T_57 = GEN_29[25:0];
  GEN_30 = {1{$random}};
  T_59 = GEN_30[2:0];
  GEN_31 = {1{$random}};
  T_61 = GEN_31[0:0];
  GEN_32 = {1{$random}};
  T_63 = GEN_32[1:0];
  GEN_33 = {1{$random}};
  T_65 = GEN_33[7:0];
  GEN_35 = {1{$random}};
  T_83 = GEN_35[0:0];
  GEN_36 = {1{$random}};
  T_85 = GEN_36[7:0];
  GEN_37 = {2{$random}};
  data_buffer_0 = GEN_37[63:0];
  GEN_46 = {2{$random}};
  data_buffer_1 = GEN_46[63:0];
  GEN_55 = {2{$random}};
  data_buffer_2 = GEN_55[63:0];
  GEN_56 = {2{$random}};
  data_buffer_3 = GEN_56[63:0];
  GEN_57 = {2{$random}};
  data_buffer_4 = GEN_57[63:0];
  GEN_58 = {2{$random}};
  data_buffer_5 = GEN_58[63:0];
  GEN_59 = {2{$random}};
  data_buffer_6 = GEN_59[63:0];
  GEN_60 = {2{$random}};
  data_buffer_7 = GEN_60[63:0];
  GEN_82 = {1{$random}};
  T_1689 = GEN_82[2:0];
  GEN_86 = {1{$random}};
  T_1733 = GEN_86[2:0];
  GEN_88 = {1{$random}};
  T_1743 = GEN_88[0:0];
  GEN_89 = {1{$random}};
  T_2166 = GEN_89[2:0];
  GEN_90 = {1{$random}};
  T_2206 = GEN_90[2:0];
  GEN_91 = {1{$random}};
  T_2216 = GEN_91[0:0];
  GEN_92 = {1{$random}};
  GEN_11 = GEN_92[25:0];
  GEN_93 = {1{$random}};
  GEN_12 = GEN_93[1:0];
  GEN_97 = {1{$random}};
  GEN_13 = GEN_97[0:0];
  GEN_99 = {1{$random}};
  GEN_14 = GEN_99[25:0];
  GEN_100 = {1{$random}};
  GEN_15 = GEN_100[2:0];
  GEN_101 = {1{$random}};
  GEN_16 = GEN_101[2:0];
  GEN_102 = {1{$random}};
  GEN_18 = GEN_102[0:0];
  GEN_105 = {1{$random}};
  GEN_19 = GEN_105[2:0];
  GEN_106 = {1{$random}};
  GEN_20 = GEN_106[11:0];
  GEN_107 = {2{$random}};
  GEN_22 = GEN_107[63:0];
  GEN_108 = {1{$random}};
  GEN_23 = GEN_108[0:0];
  GEN_109 = {1{$random}};
  GEN_24 = GEN_109[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_55 <= 4'h0;
    end else begin
      if(T_2335) begin
        T_55 <= 4'h0;
      end else begin
        if(T_1760) begin
          T_55 <= 4'h7;
        end
      end
    end
    if(reset) begin
      T_57 <= 26'h0;
    end else begin
      if(T_1760) begin
        T_57 <= io_inner_release_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1618) begin
        if(io_alloc_irel_should) begin
          T_59 <= io_inner_release_bits_r_type;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1618) begin
        if(io_alloc_irel_should) begin
          T_61 <= io_inner_release_bits_client_id;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1618) begin
        if(io_alloc_irel_should) begin
          T_63 <= io_inner_release_bits_client_xact_id;
        end
      end
    end
    if(reset) begin
      T_65 <= 8'h0;
    end else begin
      if(T_1618) begin
        if(T_1835) begin
          T_65 <= T_1860;
        end else begin
          if(io_alloc_irel_should) begin
            if(T_1800) begin
              T_65 <= T_1825;
            end else begin
              T_65 <= {{7'd0}, 1'h0};
            end
          end
        end
      end
    end
    if(reset) begin
      T_83 <= 1'h0;
    end else begin
      if(T_2087) begin
        T_83 <= 1'h0;
      end else begin
        if(T_1760) begin
          T_83 <= 1'h1;
        end
      end
    end
    if(reset) begin
      T_85 <= 8'h0;
    end else begin
      if(T_2086) begin
        T_85 <= T_2137;
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1642_0;
    end else begin
      if(T_1618) begin
        if(GEN_83 == io_inner_release_bits_addr_beat) begin
          data_buffer_0 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1642_1;
    end else begin
      if(T_1618) begin
        if(GEN_77 == io_inner_release_bits_addr_beat) begin
          data_buffer_1 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1642_2;
    end else begin
      if(T_1618) begin
        if(GEN_94 == io_inner_release_bits_addr_beat) begin
          data_buffer_2 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1642_3;
    end else begin
      if(T_1618) begin
        if(GEN_95 == io_inner_release_bits_addr_beat) begin
          data_buffer_3 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1642_4;
    end else begin
      if(T_1618) begin
        if(3'h4 == io_inner_release_bits_addr_beat) begin
          data_buffer_4 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1642_5;
    end else begin
      if(T_1618) begin
        if(3'h5 == io_inner_release_bits_addr_beat) begin
          data_buffer_5 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1642_6;
    end else begin
      if(T_1618) begin
        if(3'h6 == io_inner_release_bits_addr_beat) begin
          data_buffer_6 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1642_7;
    end else begin
      if(T_1618) begin
        if(3'h7 == io_inner_release_bits_addr_beat) begin
          data_buffer_7 <= GEN_0;
        end
      end
    end
    if(reset) begin
      T_1689 <= 3'h0;
    end else begin
      if(T_1687) begin
        T_1689 <= T_1694;
      end
    end
    if(reset) begin
      T_1733 <= 3'h0;
    end else begin
      if(T_1731) begin
        T_1733 <= T_1738;
      end
    end
    if(reset) begin
      T_1743 <= 1'h0;
    end else begin
      if(T_1752) begin
        T_1743 <= T_1755;
      end else begin
        if(T_1746) begin
          T_1743 <= T_1749;
        end
      end
    end
    if(reset) begin
      T_2166 <= 3'h0;
    end else begin
      if(T_2164) begin
        T_2166 <= T_2171;
      end
    end
    if(reset) begin
      T_2206 <= 3'h0;
    end else begin
      if(T_2204) begin
        T_2206 <= T_2211;
      end
    end
    if(reset) begin
      T_2216 <= 1'h0;
    end else begin
      if(T_2225) begin
        T_2216 <= T_2228;
      end else begin
        if(T_2219) begin
          T_2216 <= T_2222;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1628) begin
          $fwrite(32'h80000002,"Assertion failed: VoluntaryReleaseTracker accepted Release that wasn't voluntary!\n    at Broadcast.scala:78 assert(!(state === s_idle && io.inner.release.fire() && io.alloc.irel.should && !io.irel().isVoluntary()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1628) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1628) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_11(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_client_id,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_client_id,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [1:0] io_count
);
  reg [1:0] ram_client_xact_id [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_client_xact_id_T_324_data;
  wire  ram_client_xact_id_T_324_addr;
  wire  ram_client_xact_id_T_324_en;
  wire [1:0] ram_client_xact_id_T_280_data;
  wire  ram_client_xact_id_T_280_addr;
  wire  ram_client_xact_id_T_280_mask;
  wire  ram_client_xact_id_T_280_en;
  reg [2:0] ram_addr_beat [0:1];
  reg [31:0] GEN_1;
  wire [2:0] ram_addr_beat_T_324_data;
  wire  ram_addr_beat_T_324_addr;
  wire  ram_addr_beat_T_324_en;
  wire [2:0] ram_addr_beat_T_280_data;
  wire  ram_addr_beat_T_280_addr;
  wire  ram_addr_beat_T_280_mask;
  wire  ram_addr_beat_T_280_en;
  reg  ram_client_id [0:1];
  reg [31:0] GEN_2;
  wire  ram_client_id_T_324_data;
  wire  ram_client_id_T_324_addr;
  wire  ram_client_id_T_324_en;
  wire  ram_client_id_T_280_data;
  wire  ram_client_id_T_280_addr;
  wire  ram_client_id_T_280_mask;
  wire  ram_client_id_T_280_en;
  reg  ram_is_builtin_type [0:1];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_324_data;
  wire  ram_is_builtin_type_T_324_addr;
  wire  ram_is_builtin_type_T_324_en;
  wire  ram_is_builtin_type_T_280_data;
  wire  ram_is_builtin_type_T_280_addr;
  wire  ram_is_builtin_type_T_280_mask;
  wire  ram_is_builtin_type_T_280_en;
  reg [2:0] ram_a_type [0:1];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_324_data;
  wire  ram_a_type_T_324_addr;
  wire  ram_a_type_T_324_en;
  wire [2:0] ram_a_type_T_280_data;
  wire  ram_a_type_T_280_addr;
  wire  ram_a_type_T_280_mask;
  wire  ram_a_type_T_280_en;
  reg  T_272;
  reg [31:0] GEN_5;
  reg  T_274;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_277;
  wire  empty;
  wire  full;
  wire  T_278;
  wire  do_enq;
  wire  T_279;
  wire  do_deq;
  wire [1:0] T_312;
  wire  T_313;
  wire  GEN_13;
  wire [1:0] T_317;
  wire  T_318;
  wire  GEN_14;
  wire  T_319;
  wire  GEN_15;
  wire  T_321;
  wire  T_323;
  wire [1:0] T_353;
  wire  ptr_diff;
  wire  T_354;
  wire [1:0] T_355;
  assign io_enq_ready = T_323;
  assign io_deq_valid = T_321;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_324_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_324_data;
  assign io_deq_bits_client_id = ram_client_id_T_324_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_324_data;
  assign io_deq_bits_a_type = ram_a_type_T_324_data;
  assign io_count = T_355;
  assign ram_client_xact_id_T_324_addr = T_274;
  assign ram_client_xact_id_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_client_xact_id_T_324_data = ram_client_xact_id[ram_client_xact_id_T_324_addr];
  `else
  assign ram_client_xact_id_T_324_data = ram_client_xact_id_T_324_addr >= 2'h2 ? $random : ram_client_xact_id[ram_client_xact_id_T_324_addr];
  `endif
  assign ram_client_xact_id_T_280_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_280_addr = T_272;
  assign ram_client_xact_id_T_280_mask = do_enq;
  assign ram_client_xact_id_T_280_en = do_enq;
  assign ram_addr_beat_T_324_addr = T_274;
  assign ram_addr_beat_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_beat_T_324_data = ram_addr_beat[ram_addr_beat_T_324_addr];
  `else
  assign ram_addr_beat_T_324_data = ram_addr_beat_T_324_addr >= 2'h2 ? $random : ram_addr_beat[ram_addr_beat_T_324_addr];
  `endif
  assign ram_addr_beat_T_280_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_280_addr = T_272;
  assign ram_addr_beat_T_280_mask = do_enq;
  assign ram_addr_beat_T_280_en = do_enq;
  assign ram_client_id_T_324_addr = T_274;
  assign ram_client_id_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_client_id_T_324_data = ram_client_id[ram_client_id_T_324_addr];
  `else
  assign ram_client_id_T_324_data = ram_client_id_T_324_addr >= 2'h2 ? $random : ram_client_id[ram_client_id_T_324_addr];
  `endif
  assign ram_client_id_T_280_data = io_enq_bits_client_id;
  assign ram_client_id_T_280_addr = T_272;
  assign ram_client_id_T_280_mask = do_enq;
  assign ram_client_id_T_280_en = do_enq;
  assign ram_is_builtin_type_T_324_addr = T_274;
  assign ram_is_builtin_type_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_is_builtin_type_T_324_data = ram_is_builtin_type[ram_is_builtin_type_T_324_addr];
  `else
  assign ram_is_builtin_type_T_324_data = ram_is_builtin_type_T_324_addr >= 2'h2 ? $random : ram_is_builtin_type[ram_is_builtin_type_T_324_addr];
  `endif
  assign ram_is_builtin_type_T_280_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_280_addr = T_272;
  assign ram_is_builtin_type_T_280_mask = do_enq;
  assign ram_is_builtin_type_T_280_en = do_enq;
  assign ram_a_type_T_324_addr = T_274;
  assign ram_a_type_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_a_type_T_324_data = ram_a_type[ram_a_type_T_324_addr];
  `else
  assign ram_a_type_T_324_data = ram_a_type_T_324_addr >= 2'h2 ? $random : ram_a_type[ram_a_type_T_324_addr];
  `endif
  assign ram_a_type_T_280_data = io_enq_bits_a_type;
  assign ram_a_type_T_280_addr = T_272;
  assign ram_a_type_T_280_mask = do_enq;
  assign ram_a_type_T_280_en = do_enq;
  assign ptr_match = T_272 == T_274;
  assign T_277 = maybe_full == 1'h0;
  assign empty = ptr_match & T_277;
  assign full = ptr_match & maybe_full;
  assign T_278 = io_enq_ready & io_enq_valid;
  assign do_enq = T_278;
  assign T_279 = io_deq_ready & io_deq_valid;
  assign do_deq = T_279;
  assign T_312 = T_272 + 1'h1;
  assign T_313 = T_312[0:0];
  assign GEN_13 = do_enq ? T_313 : T_272;
  assign T_317 = T_274 + 1'h1;
  assign T_318 = T_317[0:0];
  assign GEN_14 = do_deq ? T_318 : T_274;
  assign T_319 = do_enq != do_deq;
  assign GEN_15 = T_319 ? do_enq : maybe_full;
  assign T_321 = empty == 1'h0;
  assign T_323 = full == 1'h0;
  assign T_353 = T_272 - T_274;
  assign ptr_diff = T_353[0:0];
  assign T_354 = maybe_full & ptr_match;
  assign T_355 = {T_354,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_0[1:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_1[2:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_client_id[initvar] = GEN_2[0:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  GEN_5 = {1{$random}};
  T_272 = GEN_5[0:0];
  GEN_6 = {1{$random}};
  T_274 = GEN_6[0:0];
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_client_xact_id_T_280_en & ram_client_xact_id_T_280_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_280_addr] <= ram_client_xact_id_T_280_data;
    end
    if(ram_addr_beat_T_280_en & ram_addr_beat_T_280_mask) begin
      ram_addr_beat[ram_addr_beat_T_280_addr] <= ram_addr_beat_T_280_data;
    end
    if(ram_client_id_T_280_en & ram_client_id_T_280_mask) begin
      ram_client_id[ram_client_id_T_280_addr] <= ram_client_id_T_280_data;
    end
    if(ram_is_builtin_type_T_280_en & ram_is_builtin_type_T_280_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_280_addr] <= ram_is_builtin_type_T_280_data;
    end
    if(ram_a_type_T_280_en & ram_a_type_T_280_mask) begin
      ram_a_type[ram_a_type_T_280_addr] <= ram_a_type_T_280_data;
    end
    if(reset) begin
      T_272 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_272 <= T_313;
      end
    end
    if(reset) begin
      T_274 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_274 <= T_318;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_319) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module BufferedBroadcastAcquireTracker(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should
);
  wire  T_44;
  reg [3:0] T_55;
  reg [31:0] GEN_30;
  reg [25:0] T_57;
  reg [31:0] GEN_31;
  reg  T_59;
  reg [31:0] GEN_39;
  reg [4:0] T_61;
  reg [31:0] GEN_40;
  reg [4:0] T_63;
  reg [31:0] GEN_41;
  reg [2:0] T_65;
  reg [31:0] GEN_45;
  reg [2:0] T_67;
  reg [31:0] GEN_59;
  wire [2:0] T_69;
  wire [1:0] T_99_client_xact_id;
  wire [2:0] T_99_addr_beat;
  wire  T_99_client_id;
  wire  T_99_is_builtin_type;
  wire [2:0] T_99_a_type;
  reg [2:0] T_129;
  reg [31:0] GEN_60;
  reg  T_131;
  reg [31:0] GEN_61;
  reg [1:0] T_133;
  reg [31:0] GEN_62;
  reg [7:0] T_135;
  reg [31:0] GEN_63;
  wire  T_144_pending;
  wire [2:0] T_144_up_idx;
  wire  T_144_up_done;
  wire [2:0] T_144_down_idx;
  wire  T_144_down_done;
  wire  T_153;
  wire [2:0] T_155;
  wire  T_157;
  wire  T_166_pending;
  wire [2:0] T_166_up_idx;
  wire  T_166_up_done;
  wire [2:0] T_166_down_idx;
  wire  T_166_down_done;
  reg [7:0] T_175;
  reg [31:0] GEN_64;
  reg [7:0] T_177;
  reg [31:0] GEN_66;
  wire  T_186_pending;
  wire [2:0] T_186_up_idx;
  wire  T_186_up_done;
  wire [2:0] T_186_down_idx;
  wire  T_186_down_done;
  reg  T_195;
  reg [31:0] GEN_67;
  reg  T_199;
  reg [31:0] GEN_68;
  reg [7:0] T_201;
  reg [31:0] GEN_70;
  wire  T_210_pending;
  wire [2:0] T_210_up_idx;
  wire  T_210_up_done;
  wire [2:0] T_210_down_idx;
  wire  T_210_down_done;
  wire [7:0] GEN_432;
  wire  T_219;
  wire  T_220;
  wire  T_221;
  wire  T_247_sharers;
  wire [1:0] T_299_state;
  wire  T_395_inner_sharers;
  wire [1:0] T_395_outer_state;
  wire  T_1733;
  wire  T_1734;
  wire  T_1735;
  wire  T_1736;
  wire [2:0] T_1745_0;
  wire  T_1747;
  wire  T_1750;
  wire  T_1751;
  wire [2:0] T_1760_0;
  wire  T_1762;
  wire  T_1765;
  wire  T_1767;
  wire [2:0] GEN_433;
  wire  T_1769;
  wire  T_1770;
  wire  T_1772;
  wire  T_1773;
  wire  T_1775;
  wire  T_1776;
  wire  T_1778;
  wire  T_1779;
  wire  T_1780;
  wire  T_1782;
  wire  T_1784;
  wire  T_1785;
  wire  T_1786;
  wire  T_1787;
  wire  T_1789;
  wire  T_1790;
  wire  T_1792;
  wire  T_1796;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [63:0] T_1817_0;
  wire [63:0] T_1817_1;
  wire [63:0] T_1817_2;
  wire [63:0] T_1817_3;
  wire [63:0] T_1817_4;
  wire [63:0] T_1817_5;
  wire [63:0] T_1817_6;
  wire [63:0] T_1817_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_71;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_72;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_73;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_74;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_78;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_79;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_80;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_81;
  wire [7:0] T_1835_0;
  wire [7:0] T_1835_1;
  wire [7:0] T_1835_2;
  wire [7:0] T_1835_3;
  wire [7:0] T_1835_4;
  wire [7:0] T_1835_5;
  wire [7:0] T_1835_6;
  wire [7:0] T_1835_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_82;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_83;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_85;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_86;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_87;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_95;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_96;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_97;
  wire  T_1841;
  wire  T_1842;
  wire  T_1844;
  wire  T_1845;
  wire  T_1847;
  wire  T_1848;
  wire  Queue_11_1_clk;
  wire  Queue_11_1_reset;
  wire  Queue_11_1_io_enq_ready;
  wire  Queue_11_1_io_enq_valid;
  wire [1:0] Queue_11_1_io_enq_bits_client_xact_id;
  wire [2:0] Queue_11_1_io_enq_bits_addr_beat;
  wire  Queue_11_1_io_enq_bits_client_id;
  wire  Queue_11_1_io_enq_bits_is_builtin_type;
  wire [2:0] Queue_11_1_io_enq_bits_a_type;
  wire  Queue_11_1_io_deq_ready;
  wire  Queue_11_1_io_deq_valid;
  wire [1:0] Queue_11_1_io_deq_bits_client_xact_id;
  wire [2:0] Queue_11_1_io_deq_bits_addr_beat;
  wire  Queue_11_1_io_deq_bits_client_id;
  wire  Queue_11_1_io_deq_bits_is_builtin_type;
  wire [2:0] Queue_11_1_io_deq_bits_a_type;
  wire [1:0] Queue_11_1_io_count;
  wire  T_1884;
  wire  T_1885;
  wire  T_1887;
  wire [2:0] T_1896_0;
  wire  T_1898;
  wire  T_1901;
  wire  T_1902;
  wire  T_1903;
  wire [7:0] T_1904;
  wire  T_1905;
  wire  T_1906;
  wire  T_1908;
  wire [2:0] T_1917_0;
  wire  T_1919;
  wire  T_1922;
  wire  T_1924;
  wire  T_1927;
  wire  T_1928;
  wire  T_1929;
  wire [1:0] T_1930_client_xact_id;
  wire [2:0] T_1930_addr_beat;
  wire  T_1930_client_id;
  wire  T_1930_is_builtin_type;
  wire [2:0] T_1930_a_type;
  wire [1:0] GEN_435;
  wire  T_1960;
  wire  T_1962;
  wire [2:0] T_1972_0;
  wire [2:0] T_1972_1;
  wire [2:0] T_1972_2;
  wire  T_1974;
  wire  T_1975;
  wire  T_1976;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire  T_1982;
  wire [7:0] GEN_436;
  wire [8:0] T_1984;
  wire [7:0] T_1985;
  wire [7:0] T_1986;
  wire [7:0] GEN_437;
  wire [7:0] T_1988;
  wire [7:0] T_1989;
  wire [7:0] T_1990;
  wire [7:0] T_1991;
  wire [2:0] T_2001_0;
  wire  T_2003;
  wire  T_2006;
  wire  T_2007;
  wire  T_2010;
  wire [7:0] T_2019;
  wire [7:0] T_2020;
  wire [7:0] GEN_32;
  wire [3:0] GEN_439;
  wire [4:0] T_2028;
  wire  T_2030;
  wire  T_2031;
  wire  T_2033;
  wire  T_2034;
  wire  T_2035;
  wire [4:0] T_2036;
  wire [4:0] T_2037;
  wire [2:0] T_2038;
  wire [2:0] T_2039;
  wire [2:0] T_2052_0;
  wire [2:0] T_2052_1;
  wire [2:0] T_2052_2;
  wire  T_2054;
  wire  T_2055;
  wire  T_2056;
  wire  T_2059;
  wire  T_2060;
  wire  T_2061;
  wire  T_2062;
  wire [7:0] GEN_440;
  wire [8:0] T_2064;
  wire [7:0] T_2065;
  wire [7:0] T_2066;
  wire [7:0] T_2070;
  wire [7:0] T_2072;
  wire [25:0] GEN_33;
  wire  GEN_34;
  wire [4:0] GEN_35;
  wire [4:0] GEN_36;
  wire [2:0] GEN_37;
  wire [2:0] GEN_38;
  wire [7:0] GEN_42;
  wire [7:0] GEN_43;
  wire [3:0] GEN_44;
  wire  T_2075;
  wire [2:0] T_2088_0;
  wire  T_2090;
  wire  T_2093;
  wire  T_2094;
  wire  T_2095;
  wire  T_2098;
  wire  T_2099;
  wire [7:0] T_2100;
  wire  skip_outer_acquire;
  wire  T_2109;
  wire [1:0] T_2110;
  wire  T_2111;
  wire [1:0] T_2112;
  wire  T_2113;
  wire [1:0] T_2114;
  wire  T_2115;
  wire [1:0] T_2116;
  wire  T_2117;
  wire [1:0] T_2118;
  wire  T_2119;
  wire [1:0] T_2120;
  wire  T_2121;
  wire [1:0] T_2122;
  wire [2:0] GEN_444;
  wire  T_2123;
  wire [1:0] T_2124;
  wire  T_2125;
  wire [1:0] T_2126;
  wire [1:0] T_2127;
  wire [25:0] T_2155_addr_block;
  wire [1:0] T_2155_p_type;
  wire  T_2155_client_id;
  wire  T_2183;
  wire [3:0] T_2184;
  wire  T_2193_pending;
  wire [2:0] T_2193_up_idx;
  wire  T_2193_up_done;
  wire [2:0] T_2193_down_idx;
  wire  T_2193_down_done;
  wire  T_2201;
  wire  T_2202;
  wire [1:0] GEN_446;
  wire [1:0] T_2204;
  wire [1:0] T_2205;
  wire [1:0] GEN_447;
  wire [1:0] T_2206;
  wire [1:0] GEN_448;
  wire [1:0] T_2207;
  wire  T_2208;
  wire  T_2211;
  reg [2:0] T_2219;
  reg [31:0] GEN_98;
  wire  T_2228;
  wire  T_2231;
  wire  T_2232;
  wire  T_2233;
  wire [2:0] T_2240_0;
  wire [2:0] T_2240_1;
  wire [2:0] T_2240_2;
  wire  T_2242;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  reg [2:0] T_2252;
  reg [31:0] GEN_99;
  wire  T_2254;
  wire [3:0] T_2256;
  wire [2:0] T_2257;
  wire [2:0] GEN_46;
  wire  T_2258;
  wire [2:0] T_2259;
  wire  T_2260;
  reg  T_2262;
  reg [31:0] GEN_100;
  wire  T_2264;
  wire  T_2265;
  wire [1:0] T_2267;
  wire  T_2268;
  wire  GEN_47;
  wire  T_2270;
  wire  T_2271;
  wire [1:0] T_2273;
  wire  T_2274;
  wire  GEN_48;
  wire  T_2276;
  wire  T_2280;
  wire  T_2282;
  wire  T_2283;
  wire [3:0] GEN_49;
  wire  T_2287;
  wire  T_2288;
  wire  T_2293;
  wire [2:0] T_2300_0;
  wire [2:0] T_2300_1;
  wire [2:0] T_2300_2;
  wire  T_2302;
  wire  T_2303;
  wire  T_2304;
  wire  T_2307;
  wire  T_2308;
  wire  T_2310;
  reg [2:0] T_2312;
  reg [31:0] GEN_101;
  wire  T_2314;
  wire [3:0] T_2316;
  wire [2:0] T_2317;
  wire [2:0] GEN_50;
  wire  T_2318;
  wire [2:0] T_2319;
  wire  T_2320;
  wire  T_2321;
  wire [3:0] GEN_452;
  wire  T_2324;
  wire  T_2325;
  wire  T_2326;
  wire  T_2327;
  wire [2:0] T_2335_0;
  wire [3:0] GEN_453;
  wire  T_2337;
  wire [1:0] T_2345_0;
  wire [1:0] T_2345_1;
  wire [3:0] GEN_454;
  wire  T_2347;
  wire [3:0] GEN_455;
  wire  T_2348;
  wire  T_2351;
  wire  T_2352;
  wire  T_2354;
  reg [2:0] T_2356;
  reg [31:0] GEN_102;
  wire  T_2358;
  wire [3:0] T_2360;
  wire [2:0] T_2361;
  wire [2:0] GEN_51;
  wire  T_2362;
  wire [2:0] T_2363;
  wire  T_2364;
  reg  T_2366;
  reg [31:0] GEN_103;
  wire  T_2368;
  wire  T_2369;
  wire [1:0] T_2371;
  wire  T_2372;
  wire  GEN_52;
  wire  T_2374;
  wire  T_2375;
  wire [1:0] T_2377;
  wire  T_2378;
  wire  GEN_53;
  wire  T_2380;
  wire  T_2382;
  wire  T_2383;
  wire [25:0] GEN_54;
  wire [3:0] GEN_55;
  wire  T_2386;
  wire [3:0] T_2392_0;
  wire [3:0] T_2392_1;
  wire  T_2394;
  wire  T_2395;
  wire  T_2398;
  wire  T_2400;
  wire  T_2401;
  wire  T_2403;
  wire  T_2404;
  wire  T_2405;
  wire  T_2407;
  wire  T_2408;
  wire  T_2411;
  wire  T_2412;
  wire  T_2414;
  wire  T_2415;
  wire [2:0] T_2422_0;
  wire [2:0] T_2422_1;
  wire [2:0] T_2422_2;
  wire  T_2424;
  wire  T_2425;
  wire  T_2426;
  wire  T_2429;
  wire  T_2430;
  wire  T_2433;
  wire  T_2435;
  wire  T_2436;
  wire  T_2437;
  wire  T_2438;
  wire [2:0] T_2445_0;
  wire [2:0] T_2445_1;
  wire [2:0] T_2445_2;
  wire  T_2447;
  wire  T_2448;
  wire  T_2449;
  wire  T_2452;
  wire  T_2453;
  wire [2:0] T_2461_0;
  wire [2:0] T_2461_1;
  wire [2:0] T_2461_2;
  wire  T_2463;
  wire  T_2464;
  wire  T_2465;
  wire  T_2468;
  wire  T_2469;
  wire  T_2470;
  wire [7:0] GEN_458;
  wire [8:0] T_2472;
  wire [7:0] T_2473;
  wire [7:0] T_2474;
  wire [7:0] T_2476;
  wire [7:0] T_2477;
  wire [7:0] T_2478;
  wire [7:0] T_2480;
  wire [2:0] GEN_56;
  wire  GEN_57;
  wire [1:0] GEN_58;
  wire [7:0] GEN_65;
  wire  T_2484;
  wire  T_2486;
  wire  T_2488;
  wire  T_2489;
  wire [2:0] T_2496_0;
  wire [2:0] T_2496_1;
  wire [2:0] T_2496_2;
  wire  T_2498;
  wire  T_2499;
  wire  T_2500;
  wire  T_2503;
  wire  T_2504;
  wire  T_2505;
  wire [7:0] GEN_460;
  wire [8:0] T_2507;
  wire [7:0] T_2508;
  wire [7:0] T_2509;
  wire [7:0] T_2513;
  wire [7:0] T_2514;
  wire [7:0] GEN_69;
  wire [2:0] GEN_75;
  wire  GEN_76;
  wire [1:0] GEN_77;
  wire [7:0] GEN_84;
  wire [3:0] T_2520_0;
  wire [3:0] T_2520_1;
  wire [3:0] T_2520_2;
  wire [3:0] T_2520_3;
  wire  T_2522;
  wire  T_2523;
  wire  T_2524;
  wire  T_2525;
  wire  T_2528;
  wire  T_2529;
  wire  T_2530;
  wire  T_2531;
  wire  T_2533;
  wire  T_2534;
  wire  T_2536;
  wire  T_2537;
  wire [2:0] T_2572_addr_beat;
  wire [25:0] T_2572_addr_block;
  wire [1:0] T_2572_client_xact_id;
  wire  T_2572_voluntary;
  wire [2:0] T_2572_r_type;
  wire [63:0] T_2572_data;
  wire  T_2572_client_id;
  wire [2:0] T_2639_addr_beat;
  wire [1:0] T_2639_client_xact_id;
  wire [2:0] T_2639_manager_xact_id;
  wire  T_2639_is_builtin_type;
  wire [3:0] T_2639_g_type;
  wire [63:0] T_2639_data;
  wire  T_2639_client_id;
  wire [3:0] T_2679_0;
  wire [3:0] T_2679_1;
  wire  T_2681;
  wire  T_2682;
  wire  T_2685;
  wire  T_2687;
  wire  T_2688;
  wire  T_2691;
  wire  T_2695;
  wire  T_2699;
  wire  T_2702;
  wire  T_2709;
  wire [2:0] T_2716_0;
  wire [2:0] T_2716_1;
  wire [2:0] T_2716_2;
  wire  T_2718;
  wire  T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [7:0] GEN_0;
  wire [7:0] GEN_88;
  wire [2:0] GEN_465;
  wire [7:0] GEN_89;
  wire [2:0] GEN_466;
  wire [7:0] GEN_90;
  wire [7:0] GEN_91;
  wire [7:0] GEN_92;
  wire [7:0] GEN_93;
  wire [7:0] GEN_94;
  wire  T_2726;
  wire [7:0] GEN_1;
  wire  T_2727;
  wire [7:0] GEN_2;
  wire  T_2728;
  wire [7:0] GEN_3;
  wire  T_2729;
  wire [7:0] GEN_4;
  wire  T_2730;
  wire [7:0] GEN_5;
  wire  T_2731;
  wire [7:0] GEN_6;
  wire  T_2732;
  wire [7:0] GEN_7;
  wire  T_2733;
  wire [7:0] GEN_488;
  wire [8:0] T_2735;
  wire [7:0] T_2736;
  wire [7:0] GEN_489;
  wire [8:0] T_2738;
  wire [7:0] T_2739;
  wire [7:0] GEN_490;
  wire [8:0] T_2741;
  wire [7:0] T_2742;
  wire [7:0] GEN_491;
  wire [8:0] T_2744;
  wire [7:0] T_2745;
  wire [7:0] GEN_492;
  wire [8:0] T_2747;
  wire [7:0] T_2748;
  wire [7:0] GEN_493;
  wire [8:0] T_2750;
  wire [7:0] T_2751;
  wire [7:0] GEN_494;
  wire [8:0] T_2753;
  wire [7:0] T_2754;
  wire [7:0] GEN_495;
  wire [8:0] T_2756;
  wire [7:0] T_2757;
  wire [7:0] T_2763_0;
  wire [7:0] T_2763_1;
  wire [7:0] T_2763_2;
  wire [7:0] T_2763_3;
  wire [7:0] T_2763_4;
  wire [7:0] T_2763_5;
  wire [7:0] T_2763_6;
  wire [7:0] T_2763_7;
  wire [15:0] T_2765;
  wire [15:0] T_2766;
  wire [31:0] T_2767;
  wire [15:0] T_2768;
  wire [15:0] T_2769;
  wire [31:0] T_2770;
  wire [63:0] T_2771;
  wire [63:0] T_2772;
  wire [63:0] T_2773;
  wire [63:0] GEN_8;
  wire [63:0] GEN_144;
  wire [63:0] GEN_145;
  wire [63:0] GEN_146;
  wire [63:0] GEN_147;
  wire [63:0] GEN_148;
  wire [63:0] GEN_149;
  wire [63:0] GEN_150;
  wire [63:0] T_2774;
  wire [63:0] T_2775;
  wire [63:0] GEN_9;
  wire [63:0] GEN_151;
  wire [63:0] GEN_152;
  wire [63:0] GEN_153;
  wire [63:0] GEN_154;
  wire [63:0] GEN_155;
  wire [63:0] GEN_156;
  wire [63:0] GEN_157;
  wire [63:0] GEN_158;
  wire [63:0] GEN_177;
  wire [63:0] GEN_178;
  wire [63:0] GEN_179;
  wire [63:0] GEN_180;
  wire [63:0] GEN_181;
  wire [63:0] GEN_182;
  wire [63:0] GEN_183;
  wire [63:0] GEN_184;
  wire [1:0] T_2806_state;
  wire  T_2832;
  wire  T_2833;
  wire [2:0] T_2839_0;
  wire [2:0] T_2839_1;
  wire [2:0] T_2839_2;
  wire  T_2841;
  wire  T_2842;
  wire  T_2843;
  wire  T_2846;
  wire  T_2847;
  wire  T_2848;
  wire [7:0] GEN_503;
  wire [8:0] T_2850;
  wire [7:0] T_2851;
  wire [7:0] T_2852;
  wire [7:0] T_2854;
  wire [7:0] T_2855;
  wire [7:0] T_2856;
  wire [7:0] T_2857;
  wire [2:0] T_2865_0;
  wire [2:0] T_2865_1;
  wire [2:0] T_2865_2;
  wire  T_2867;
  wire  T_2868;
  wire  T_2869;
  wire  T_2872;
  wire  T_2873;
  wire  T_2874;
  wire [7:0] GEN_505;
  wire [8:0] T_2877;
  wire [7:0] T_2878;
  wire [7:0] T_2881;
  wire [7:0] T_2882;
  wire [7:0] T_2883;
  wire [7:0] GEN_191;
  wire  GEN_193;
  wire  T_2893;
  wire [2:0] T_2900_0;
  wire [2:0] T_2900_1;
  wire [2:0] T_2900_2;
  wire  T_2902;
  wire  T_2903;
  wire  T_2904;
  wire  T_2907;
  wire  T_2908;
  wire  T_2910;
  reg [2:0] T_2912;
  reg [31:0] GEN_104;
  wire  T_2914;
  wire [3:0] T_2916;
  wire [2:0] T_2917;
  wire [2:0] GEN_194;
  wire  T_2918;
  wire [2:0] T_2919;
  wire  T_2920;
  wire  T_2923;
  wire  T_2924;
  wire  T_2925;
  wire [2:0] T_2933_0;
  wire [3:0] GEN_510;
  wire  T_2935;
  wire  T_2943_0;
  wire [3:0] GEN_511;
  wire  T_2945;
  wire  T_2948;
  wire  T_2950;
  reg [2:0] T_2952;
  reg [31:0] GEN_105;
  wire  T_2954;
  wire [3:0] T_2956;
  wire [2:0] T_2957;
  wire [2:0] GEN_195;
  wire  T_2958;
  wire [2:0] T_2959;
  wire  T_2960;
  reg  T_2962;
  reg [31:0] GEN_106;
  wire  T_2964;
  wire  T_2965;
  wire [1:0] T_2967;
  wire  T_2968;
  wire  GEN_196;
  wire  T_2970;
  wire  T_2971;
  wire [1:0] T_2973;
  wire  T_2974;
  wire  GEN_197;
  wire  T_2976;
  wire  T_2977;
  wire [2:0] T_2983_0;
  wire [2:0] T_2983_1;
  wire [2:0] T_2983_2;
  wire  T_2985;
  wire  T_2986;
  wire  T_2987;
  wire  T_2990;
  wire  T_2991;
  wire [7:0] T_2992;
  wire  T_2993;
  wire  T_2995;
  wire  T_2996;
  wire [1:0] T_3004_0;
  wire  T_3006;
  wire [2:0] T_3009;
  wire [2:0] T_3045_addr_beat;
  wire [25:0] T_3045_addr_block;
  wire [2:0] T_3045_client_xact_id;
  wire  T_3045_voluntary;
  wire [2:0] T_3045_r_type;
  wire [63:0] T_3045_data;
  wire [63:0] GEN_10;
  wire [63:0] GEN_198;
  wire [63:0] GEN_199;
  wire [63:0] GEN_200;
  wire [63:0] GEN_201;
  wire [63:0] GEN_202;
  wire [63:0] GEN_203;
  wire [63:0] GEN_204;
  wire  T_3074;
  wire  T_3076;
  wire [2:0] T_3087_0;
  wire  T_3089;
  wire  T_3092;
  wire  T_3093;
  reg [2:0] T_3095;
  reg [31:0] GEN_107;
  wire  T_3097;
  wire [3:0] T_3099;
  wire [2:0] T_3100;
  wire [2:0] GEN_205;
  wire  T_3101;
  wire [2:0] T_3102;
  wire  T_3103;
  wire  T_3109;
  wire  T_3110;
  wire [2:0] T_3118_0;
  wire [3:0] GEN_518;
  wire  T_3120;
  wire  T_3128_0;
  wire [3:0] GEN_519;
  wire  T_3130;
  wire  T_3133;
  wire  T_3135;
  reg [2:0] T_3137;
  reg [31:0] GEN_108;
  wire  T_3139;
  wire [3:0] T_3141;
  wire [2:0] T_3142;
  wire [2:0] GEN_206;
  wire  T_3143;
  wire [2:0] T_3144;
  wire  T_3145;
  reg  T_3147;
  reg [31:0] GEN_109;
  wire  T_3149;
  wire  T_3150;
  wire [1:0] T_3152;
  wire  T_3153;
  wire  GEN_207;
  wire  T_3155;
  wire  T_3156;
  wire [1:0] T_3158;
  wire  T_3159;
  wire  GEN_208;
  wire  T_3161;
  wire  T_3162;
  wire [7:0] T_3163;
  wire  T_3164;
  wire  T_3166;
  wire  T_3168;
  wire  T_3169;
  wire  T_3172;
  wire  T_3173;
  wire  T_3174;
  wire  T_3175;
  wire  T_3176;
  wire  T_3177;
  wire  T_3178;
  wire  T_3179;
  wire  T_3180;
  wire  T_3181;
  wire  T_3182;
  wire [5:0] T_3185;
  wire [25:0] T_3216_addr_block;
  wire [2:0] T_3216_client_xact_id;
  wire [2:0] T_3216_addr_beat;
  wire  T_3216_is_builtin_type;
  wire [2:0] T_3216_a_type;
  wire [11:0] T_3216_union;
  wire [63:0] T_3216_data;
  wire [7:0] GEN_11;
  wire [7:0] GEN_209;
  wire [7:0] GEN_210;
  wire [7:0] GEN_211;
  wire [7:0] GEN_212;
  wire [7:0] GEN_213;
  wire [7:0] GEN_214;
  wire [7:0] GEN_215;
  wire [5:0] T_3281;
  wire [5:0] T_3282;
  wire [11:0] T_3283;
  wire [7:0] T_3285;
  wire [8:0] T_3286;
  wire [8:0] T_3288;
  wire [5:0] T_3300;
  wire [5:0] T_3302;
  wire [11:0] T_3304;
  wire [11:0] T_3306;
  wire [11:0] T_3308;
  wire [11:0] T_3310;
  wire [11:0] T_3312;
  wire [25:0] T_3341_addr_block;
  wire [2:0] T_3341_client_xact_id;
  wire [2:0] T_3341_addr_beat;
  wire  T_3341_is_builtin_type;
  wire [2:0] T_3341_a_type;
  wire [11:0] T_3341_union;
  wire [63:0] T_3341_data;
  wire [63:0] GEN_12;
  wire [63:0] GEN_216;
  wire [63:0] GEN_217;
  wire [63:0] GEN_218;
  wire [63:0] GEN_219;
  wire [63:0] GEN_220;
  wire [63:0] GEN_221;
  wire [63:0] GEN_222;
  wire [25:0] T_3369_addr_block;
  wire [2:0] T_3369_client_xact_id;
  wire [2:0] T_3369_addr_beat;
  wire  T_3369_is_builtin_type;
  wire [2:0] T_3369_a_type;
  wire [11:0] T_3369_union;
  wire [63:0] T_3369_data;
  wire  T_3398;
  wire [3:0] GEN_223;
  wire [2:0] T_3408_0;
  wire [2:0] T_3408_1;
  wire [3:0] GEN_527;
  wire  T_3410;
  wire [3:0] GEN_528;
  wire  T_3411;
  wire  T_3414;
  wire  T_3420_0;
  wire [3:0] GEN_529;
  wire  T_3422;
  wire  T_3425;
  wire  T_3426;
  wire [7:0] GEN_13;
  wire [7:0] GEN_224;
  wire [7:0] GEN_225;
  wire [7:0] GEN_226;
  wire [7:0] GEN_227;
  wire [7:0] GEN_228;
  wire [7:0] GEN_229;
  wire [7:0] GEN_230;
  wire  T_3427;
  wire [7:0] GEN_14;
  wire  T_3428;
  wire [7:0] GEN_15;
  wire  T_3429;
  wire [7:0] GEN_16;
  wire  T_3430;
  wire [7:0] GEN_17;
  wire  T_3431;
  wire [7:0] GEN_18;
  wire  T_3432;
  wire [7:0] GEN_19;
  wire  T_3433;
  wire [7:0] GEN_20;
  wire  T_3434;
  wire [7:0] GEN_554;
  wire [8:0] T_3436;
  wire [7:0] T_3437;
  wire [7:0] GEN_555;
  wire [8:0] T_3439;
  wire [7:0] T_3440;
  wire [7:0] GEN_556;
  wire [8:0] T_3442;
  wire [7:0] T_3443;
  wire [7:0] GEN_557;
  wire [8:0] T_3445;
  wire [7:0] T_3446;
  wire [7:0] GEN_558;
  wire [8:0] T_3448;
  wire [7:0] T_3449;
  wire [7:0] GEN_559;
  wire [8:0] T_3451;
  wire [7:0] T_3452;
  wire [7:0] GEN_560;
  wire [8:0] T_3454;
  wire [7:0] T_3455;
  wire [7:0] GEN_561;
  wire [8:0] T_3457;
  wire [7:0] T_3458;
  wire [7:0] T_3464_0;
  wire [7:0] T_3464_1;
  wire [7:0] T_3464_2;
  wire [7:0] T_3464_3;
  wire [7:0] T_3464_4;
  wire [7:0] T_3464_5;
  wire [7:0] T_3464_6;
  wire [7:0] T_3464_7;
  wire [15:0] T_3466;
  wire [15:0] T_3467;
  wire [31:0] T_3468;
  wire [15:0] T_3469;
  wire [15:0] T_3470;
  wire [31:0] T_3471;
  wire [63:0] T_3472;
  wire [63:0] T_3473;
  wire [63:0] T_3474;
  wire [63:0] GEN_21;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [63:0] GEN_286;
  wire [63:0] T_3475;
  wire [63:0] T_3476;
  wire [63:0] GEN_22;
  wire [63:0] GEN_287;
  wire [63:0] GEN_288;
  wire [63:0] GEN_289;
  wire [63:0] GEN_290;
  wire [63:0] GEN_291;
  wire [63:0] GEN_292;
  wire [63:0] GEN_293;
  wire [63:0] GEN_294;
  wire [63:0] GEN_313;
  wire [63:0] GEN_314;
  wire [63:0] GEN_315;
  wire [63:0] GEN_316;
  wire [63:0] GEN_317;
  wire [63:0] GEN_318;
  wire [63:0] GEN_319;
  wire [63:0] GEN_320;
  wire  T_3477;
  wire  T_3478;
  wire  T_3489;
  wire  T_3491;
  wire [2:0] T_3499_0;
  wire [3:0] GEN_570;
  wire  T_3501;
  wire [1:0] T_3509_0;
  wire [1:0] T_3509_1;
  wire [3:0] GEN_571;
  wire  T_3511;
  wire [3:0] GEN_572;
  wire  T_3512;
  wire  T_3515;
  wire  T_3516;
  wire  T_3518;
  reg [2:0] T_3520;
  reg [31:0] GEN_110;
  wire  T_3522;
  wire [3:0] T_3524;
  wire [2:0] T_3525;
  wire [2:0] GEN_321;
  wire  T_3526;
  wire [2:0] T_3527;
  wire  T_3528;
  wire  T_3529;
  reg [2:0] T_3535;
  reg [31:0] GEN_111;
  reg  T_3545;
  reg [31:0] GEN_112;
  wire  T_3547;
  wire  T_3548;
  wire [1:0] T_3550;
  wire  T_3551;
  wire  GEN_323;
  wire  T_3553;
  wire  T_3554;
  wire [1:0] T_3556;
  wire  T_3557;
  wire  GEN_324;
  wire  T_3559;
  wire  T_3564;
  wire [2:0] T_3573_0;
  wire [2:0] T_3573_1;
  wire [3:0] GEN_575;
  wire  T_3575;
  wire [3:0] GEN_576;
  wire  T_3576;
  wire  T_3579;
  wire [1:0] T_3585_0;
  wire [1:0] T_3585_1;
  wire [3:0] GEN_577;
  wire  T_3587;
  wire [3:0] GEN_578;
  wire  T_3588;
  wire  T_3591;
  wire  T_3592;
  wire  T_3593;
  wire [7:0] GEN_579;
  wire [8:0] T_3595;
  wire [7:0] T_3596;
  wire [7:0] T_3597;
  wire [7:0] T_3599;
  wire [7:0] T_3600;
  wire [7:0] T_3601;
  wire [7:0] T_3602;
  wire [2:0] T_3610_0;
  wire [2:0] T_3610_1;
  wire [2:0] T_3610_2;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3617;
  wire  T_3618;
  wire  T_3619;
  wire [7:0] GEN_581;
  wire [8:0] T_3622;
  wire [7:0] T_3623;
  wire [7:0] T_3626;
  wire [7:0] T_3627;
  wire [2:0] T_3637_0;
  wire [2:0] T_3637_1;
  wire [3:0] GEN_583;
  wire  T_3639;
  wire [3:0] GEN_584;
  wire  T_3640;
  wire  T_3643;
  wire  T_3649_0;
  wire [3:0] GEN_585;
  wire  T_3651;
  wire  T_3654;
  wire  T_3655;
  wire [7:0] GEN_586;
  wire [8:0] T_3658;
  wire [7:0] T_3659;
  wire [7:0] T_3661;
  wire [7:0] T_3662;
  wire [7:0] T_3663;
  wire [7:0] T_3664;
  wire [7:0] GEN_335;
  wire  T_3666;
  wire  T_3667;
  wire  T_3670;
  wire  T_3672;
  wire  T_3689;
  wire [2:0] T_3690;
  wire  T_3691;
  wire [2:0] T_3692;
  wire  T_3693;
  wire [2:0] T_3694;
  wire  T_3695;
  wire [2:0] T_3696;
  wire  T_3697;
  wire [2:0] T_3698;
  wire  T_3699;
  wire [2:0] T_3700;
  wire  T_3701;
  wire [2:0] T_3702;
  wire  T_3703;
  wire [1:0] T_3708;
  wire [2:0] T_3709;
  wire [2:0] T_3741_addr_beat;
  wire [1:0] T_3741_client_xact_id;
  wire [2:0] T_3741_manager_xact_id;
  wire  T_3741_is_builtin_type;
  wire [3:0] T_3741_g_type;
  wire [63:0] T_3741_data;
  wire  T_3741_client_id;
  wire [63:0] GEN_23;
  wire [63:0] GEN_336;
  wire [63:0] GEN_337;
  wire [63:0] GEN_338;
  wire [63:0] GEN_339;
  wire [63:0] GEN_340;
  wire [63:0] GEN_341;
  wire [63:0] GEN_342;
  wire [2:0] T_3780_0;
  wire [3:0] GEN_594;
  wire  T_3782;
  wire [1:0] T_3790_0;
  wire [1:0] T_3790_1;
  wire [3:0] GEN_595;
  wire  T_3792;
  wire [3:0] GEN_596;
  wire  T_3793;
  wire  T_3796;
  wire  T_3797;
  wire  T_3799;
  reg [2:0] T_3801;
  reg [31:0] GEN_113;
  wire  T_3803;
  wire [3:0] T_3805;
  wire [2:0] T_3806;
  wire [2:0] GEN_343;
  wire  T_3807;
  wire [2:0] T_3808;
  wire  T_3809;
  wire  T_3814;
  wire  T_3816;
  wire [2:0] T_3824_0;
  wire [2:0] T_3824_1;
  wire [3:0] GEN_598;
  wire  T_3826;
  wire [3:0] GEN_599;
  wire  T_3827;
  wire  T_3830;
  wire [1:0] T_3836_0;
  wire [1:0] T_3836_1;
  wire [3:0] GEN_600;
  wire  T_3838;
  wire [3:0] GEN_601;
  wire  T_3839;
  wire  T_3842;
  wire  T_3843;
  wire [7:0] T_3844;
  wire  T_3845;
  wire  T_3846;
  wire  T_3847;
  wire  GEN_348;
  wire  GEN_349;
  wire [2:0] GEN_350;
  wire [1:0] GEN_351;
  wire [2:0] GEN_352;
  wire  GEN_353;
  wire [3:0] GEN_354;
  wire [63:0] GEN_355;
  wire  GEN_356;
  wire  GEN_361;
  wire  T_3854;
  wire [1:0] GEN_362;
  wire [2:0] T_3869_0;
  wire  T_3871;
  wire  T_3874;
  wire  T_3875;
  wire  T_3876;
  wire  T_3879;
  wire  T_3881;
  wire  T_3882;
  wire [2:0] T_3892_0;
  wire [2:0] T_3892_1;
  wire [2:0] T_3892_2;
  wire  T_3894;
  wire  T_3895;
  wire  T_3896;
  wire  T_3899;
  wire  T_3900;
  wire  T_3901;
  wire  T_3902;
  wire  T_3903;
  wire  T_3905;
  wire  T_3906;
  wire [8:0] T_3910;
  wire [7:0] T_3911;
  wire [7:0] T_3917_0;
  wire  T_3925;
  wire [7:0] T_3926;
  wire [7:0] T_3928;
  wire [7:0] T_3929;
  wire  T_3930;
  wire  T_3931;
  wire  T_3932;
  wire  T_3933;
  wire  T_3934;
  wire  T_3935;
  wire  T_3936;
  wire  T_3937;
  wire [7:0] GEN_603;
  wire [8:0] T_3939;
  wire [7:0] T_3940;
  wire [7:0] GEN_604;
  wire [8:0] T_3942;
  wire [7:0] T_3943;
  wire [7:0] GEN_605;
  wire [8:0] T_3945;
  wire [7:0] T_3946;
  wire [7:0] GEN_606;
  wire [8:0] T_3948;
  wire [7:0] T_3949;
  wire [7:0] GEN_607;
  wire [8:0] T_3951;
  wire [7:0] T_3952;
  wire [7:0] GEN_608;
  wire [8:0] T_3954;
  wire [7:0] T_3955;
  wire [7:0] GEN_609;
  wire [8:0] T_3957;
  wire [7:0] T_3958;
  wire [7:0] GEN_610;
  wire [8:0] T_3960;
  wire [7:0] T_3961;
  wire [7:0] T_3967_0;
  wire [7:0] T_3967_1;
  wire [7:0] T_3967_2;
  wire [7:0] T_3967_3;
  wire [7:0] T_3967_4;
  wire [7:0] T_3967_5;
  wire [7:0] T_3967_6;
  wire [7:0] T_3967_7;
  wire [15:0] T_3969;
  wire [15:0] T_3970;
  wire [31:0] T_3971;
  wire [15:0] T_3972;
  wire [15:0] T_3973;
  wire [31:0] T_3974;
  wire [63:0] T_3975;
  wire [63:0] T_3976;
  wire [63:0] GEN_24;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [63:0] GEN_366;
  wire [63:0] GEN_367;
  wire [63:0] GEN_368;
  wire [63:0] GEN_369;
  wire [63:0] T_3977;
  wire [63:0] T_3978;
  wire [63:0] T_3979;
  wire [63:0] GEN_25;
  wire [63:0] GEN_370;
  wire [63:0] GEN_371;
  wire [63:0] GEN_372;
  wire [63:0] GEN_373;
  wire [63:0] GEN_374;
  wire [63:0] GEN_375;
  wire [63:0] GEN_376;
  wire [63:0] GEN_377;
  wire [7:0] T_3993_0;
  wire [7:0] T_4005;
  wire [7:0] GEN_26;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [7:0] GEN_381;
  wire [7:0] GEN_382;
  wire [7:0] GEN_383;
  wire [7:0] GEN_384;
  wire [7:0] T_4006;
  wire [7:0] GEN_27;
  wire [7:0] GEN_385;
  wire [7:0] GEN_386;
  wire [7:0] GEN_387;
  wire [7:0] GEN_388;
  wire [7:0] GEN_389;
  wire [7:0] GEN_390;
  wire [7:0] GEN_391;
  wire [7:0] GEN_392;
  wire [63:0] GEN_404;
  wire [63:0] GEN_405;
  wire [63:0] GEN_406;
  wire [63:0] GEN_407;
  wire [63:0] GEN_408;
  wire [63:0] GEN_409;
  wire [63:0] GEN_410;
  wire [63:0] GEN_411;
  wire [7:0] GEN_415;
  wire [7:0] GEN_416;
  wire [7:0] GEN_417;
  wire [7:0] GEN_418;
  wire [7:0] GEN_419;
  wire [7:0] GEN_420;
  wire [7:0] GEN_421;
  wire [7:0] GEN_422;
  wire  T_4009;
  wire  T_4010;
  wire  T_4011;
  wire  T_4012;
  wire  T_4013;
  wire  T_4014;
  wire  T_4015;
  wire  T_4017;
  wire  T_4019;
  wire [3:0] GEN_423;
  wire [7:0] GEN_424;
  wire [7:0] GEN_425;
  wire [7:0] GEN_426;
  wire [7:0] GEN_427;
  wire [7:0] GEN_428;
  wire [7:0] GEN_429;
  wire [7:0] GEN_430;
  wire [7:0] GEN_431;
  reg  GEN_28;
  reg [31:0] GEN_114;
  reg  GEN_29;
  reg [31:0] GEN_115;
  Queue_11 Queue_11_1 (
    .clk(Queue_11_1_clk),
    .reset(Queue_11_1_reset),
    .io_enq_ready(Queue_11_1_io_enq_ready),
    .io_enq_valid(Queue_11_1_io_enq_valid),
    .io_enq_bits_client_xact_id(Queue_11_1_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(Queue_11_1_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(Queue_11_1_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(Queue_11_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(Queue_11_1_io_enq_bits_a_type),
    .io_deq_ready(Queue_11_1_io_deq_ready),
    .io_deq_valid(Queue_11_1_io_deq_valid),
    .io_deq_bits_client_xact_id(Queue_11_1_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(Queue_11_1_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(Queue_11_1_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(Queue_11_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(Queue_11_1_io_deq_bits_a_type),
    .io_count(Queue_11_1_io_count)
  );
  assign io_inner_acquire_ready = T_2099;
  assign io_inner_grant_valid = GEN_361;
  assign io_inner_grant_bits_addr_beat = GEN_350;
  assign io_inner_grant_bits_client_xact_id = GEN_351;
  assign io_inner_grant_bits_manager_xact_id = GEN_352;
  assign io_inner_grant_bits_is_builtin_type = GEN_353;
  assign io_inner_grant_bits_g_type = GEN_354;
  assign io_inner_grant_bits_data = GEN_355;
  assign io_inner_grant_bits_client_id = GEN_356;
  assign io_inner_finish_ready = T_2977;
  assign io_inner_probe_valid = T_2211;
  assign io_inner_probe_bits_addr_block = T_2155_addr_block;
  assign io_inner_probe_bits_p_type = T_2155_p_type;
  assign io_inner_probe_bits_client_id = T_2155_client_id;
  assign io_inner_release_ready = T_2709;
  assign io_outer_acquire_valid = T_3169;
  assign io_outer_acquire_bits_addr_block = T_3369_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3369_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3369_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3369_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3369_a_type;
  assign io_outer_acquire_bits_union = T_3369_union;
  assign io_outer_acquire_bits_data = T_3369_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2996;
  assign io_outer_release_bits_addr_beat = T_3045_addr_beat;
  assign io_outer_release_bits_addr_block = T_3045_addr_block;
  assign io_outer_release_bits_client_xact_id = T_3045_client_xact_id;
  assign io_outer_release_bits_voluntary = T_3045_voluntary;
  assign io_outer_release_bits_r_type = T_3045_r_type;
  assign io_outer_release_bits_data = T_3045_data;
  assign io_outer_grant_ready = T_2977;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_28;
  assign io_outer_finish_bits_manager_id = GEN_29;
  assign io_alloc_iacq_matches = T_1842;
  assign io_alloc_iacq_can = T_1733;
  assign io_alloc_irel_matches = T_1845;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1848;
  assign io_alloc_oprb_can = 1'h0;
  assign T_44 = T_4017;
  assign T_69 = T_99_addr_beat;
  assign T_99_client_xact_id = T_1930_client_xact_id;
  assign T_99_addr_beat = T_1930_addr_beat;
  assign T_99_client_id = T_1930_client_id;
  assign T_99_is_builtin_type = T_1930_is_builtin_type;
  assign T_99_a_type = T_1930_a_type;
  assign T_144_pending = T_2380;
  assign T_144_up_idx = T_2319;
  assign T_144_up_done = T_2320;
  assign T_144_down_idx = T_2363;
  assign T_144_down_done = T_2364;
  assign T_153 = T_1960;
  assign T_155 = T_3808;
  assign T_157 = T_3809;
  assign T_166_pending = T_3559;
  assign T_166_up_idx = T_3527;
  assign T_166_up_done = T_3528;
  assign T_166_down_idx = 3'h0;
  assign T_166_down_done = T_3529;
  assign T_186_pending = T_3161;
  assign T_186_up_idx = T_3102;
  assign T_186_up_done = T_3103;
  assign T_186_down_idx = T_3144;
  assign T_186_down_done = T_3145;
  assign T_210_pending = T_2976;
  assign T_210_up_idx = T_2919;
  assign T_210_up_done = T_2920;
  assign T_210_down_idx = T_2959;
  assign T_210_down_done = T_2960;
  assign GEN_432 = {{7'd0}, 1'h0};
  assign T_219 = T_201 != GEN_432;
  assign T_220 = T_199 | T_219;
  assign T_221 = T_220 | T_210_pending;
  assign T_247_sharers = 1'h0;
  assign T_299_state = {{1'd0}, 1'h0};
  assign T_395_inner_sharers = T_247_sharers;
  assign T_395_outer_state = T_299_state;
  assign T_1733 = T_55 == 4'h0;
  assign T_1734 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1735 = T_1733 & T_1734;
  assign T_1736 = T_1735 & io_alloc_iacq_should;
  assign T_1745_0 = 3'h3;
  assign T_1747 = T_1745_0 == io_inner_acquire_bits_a_type;
  assign T_1750 = io_inner_acquire_bits_is_builtin_type & T_1747;
  assign T_1751 = T_1736 & T_1750;
  assign T_1760_0 = 3'h3;
  assign T_1762 = T_1760_0 == io_inner_acquire_bits_a_type;
  assign T_1765 = io_inner_acquire_bits_is_builtin_type & T_1762;
  assign T_1767 = T_1765 == 1'h0;
  assign GEN_433 = {{2'd0}, 1'h0};
  assign T_1769 = io_inner_acquire_bits_addr_beat == GEN_433;
  assign T_1770 = T_1767 | T_1769;
  assign T_1772 = T_1770 == 1'h0;
  assign T_1773 = T_1751 & T_1772;
  assign T_1775 = T_1773 == 1'h0;
  assign T_1776 = T_1775 | reset;
  assign T_1778 = T_1776 == 1'h0;
  assign T_1779 = T_55 != 4'h0;
  assign T_1780 = T_1779 & T_153;
  assign T_1782 = T_99_a_type == 3'h5;
  assign T_1784 = T_99_a_type == 3'h6;
  assign T_1785 = T_1782 | T_1784;
  assign T_1786 = T_99_is_builtin_type & T_1785;
  assign T_1787 = T_1780 & T_1786;
  assign T_1789 = T_1787 == 1'h0;
  assign T_1790 = T_1789 | reset;
  assign T_1792 = T_1790 == 1'h0;
  assign T_1796 = T_99_a_type == 3'h4;
  assign T_1797 = T_99_is_builtin_type & T_1796;
  assign T_1798 = T_1780 & T_1797;
  assign T_1800 = T_1798 == 1'h0;
  assign T_1801 = T_1800 | reset;
  assign T_1803 = T_1801 == 1'h0;
  assign T_1817_0 = 64'h0;
  assign T_1817_1 = 64'h0;
  assign T_1817_2 = 64'h0;
  assign T_1817_3 = 64'h0;
  assign T_1817_4 = 64'h0;
  assign T_1817_5 = 64'h0;
  assign T_1817_6 = 64'h0;
  assign T_1817_7 = 64'h0;
  assign T_1835_0 = 8'h0;
  assign T_1835_1 = 8'h0;
  assign T_1835_2 = 8'h0;
  assign T_1835_3 = 8'h0;
  assign T_1835_4 = 8'h0;
  assign T_1835_5 = 8'h0;
  assign T_1835_6 = 8'h0;
  assign T_1835_7 = 8'h0;
  assign T_1841 = io_inner_acquire_bits_addr_block == T_57;
  assign T_1842 = T_1779 & T_1841;
  assign T_1844 = io_inner_release_bits_addr_block == T_57;
  assign T_1845 = T_1779 & T_1844;
  assign T_1847 = io_outer_probe_bits_addr_block == T_57;
  assign T_1848 = T_1779 & T_1847;
  assign Queue_11_1_clk = clk;
  assign Queue_11_1_reset = reset;
  assign Queue_11_1_io_enq_valid = T_1929;
  assign Queue_11_1_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign Queue_11_1_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign Queue_11_1_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign Queue_11_1_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign Queue_11_1_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign Queue_11_1_io_deq_ready = GEN_349;
  assign T_1884 = T_1733 & io_alloc_iacq_should;
  assign T_1885 = T_1884 & io_inner_acquire_valid;
  assign T_1887 = T_99_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1896_0 = 3'h3;
  assign T_1898 = T_1896_0 == T_99_a_type;
  assign T_1901 = T_99_is_builtin_type & T_1898;
  assign T_1902 = T_1887 & T_1901;
  assign T_1903 = T_1902 & T_153;
  assign T_1904 = T_175 >> io_inner_acquire_bits_addr_beat;
  assign T_1905 = T_1904[0];
  assign T_1906 = T_1903 & T_1905;
  assign T_1908 = T_1906 & io_inner_acquire_valid;
  assign T_1917_0 = 3'h3;
  assign T_1919 = T_1917_0 == io_inner_acquire_bits_a_type;
  assign T_1922 = io_inner_acquire_bits_is_builtin_type & T_1919;
  assign T_1924 = T_1922 == 1'h0;
  assign T_1927 = T_1924 | T_1769;
  assign T_1928 = T_1908 & T_1927;
  assign T_1929 = T_1885 | T_1928;
  assign T_1930_client_xact_id = Queue_11_1_io_deq_valid ? Queue_11_1_io_deq_bits_client_xact_id : Queue_11_1_io_enq_bits_client_xact_id;
  assign T_1930_addr_beat = Queue_11_1_io_deq_valid ? Queue_11_1_io_deq_bits_addr_beat : Queue_11_1_io_enq_bits_addr_beat;
  assign T_1930_client_id = Queue_11_1_io_deq_valid ? Queue_11_1_io_deq_bits_client_id : Queue_11_1_io_enq_bits_client_id;
  assign T_1930_is_builtin_type = Queue_11_1_io_deq_valid ? Queue_11_1_io_deq_bits_is_builtin_type : Queue_11_1_io_enq_bits_is_builtin_type;
  assign T_1930_a_type = Queue_11_1_io_deq_valid ? Queue_11_1_io_deq_bits_a_type : Queue_11_1_io_enq_bits_a_type;
  assign GEN_435 = {{1'd0}, 1'h0};
  assign T_1960 = Queue_11_1_io_count > GEN_435;
  assign T_1962 = T_1779 | io_alloc_iacq_should;
  assign T_1972_0 = 3'h2;
  assign T_1972_1 = 3'h3;
  assign T_1972_2 = 3'h4;
  assign T_1974 = T_1972_0 == io_inner_acquire_bits_a_type;
  assign T_1975 = T_1972_1 == io_inner_acquire_bits_a_type;
  assign T_1976 = T_1972_2 == io_inner_acquire_bits_a_type;
  assign T_1979 = T_1974 | T_1975;
  assign T_1980 = T_1979 | T_1976;
  assign T_1981 = io_inner_acquire_bits_is_builtin_type & T_1980;
  assign T_1982 = T_1734 & T_1981;
  assign GEN_436 = {{7'd0}, T_1982};
  assign T_1984 = 8'h0 - GEN_436;
  assign T_1985 = T_1984[7:0];
  assign T_1986 = ~ T_1985;
  assign GEN_437 = {{7'd0}, 1'h1};
  assign T_1988 = GEN_437 << io_inner_acquire_bits_addr_beat;
  assign T_1989 = ~ T_1988;
  assign T_1990 = T_1986 | T_1989;
  assign T_1991 = T_175 & T_1990;
  assign T_2001_0 = 3'h3;
  assign T_2003 = T_2001_0 == io_inner_acquire_bits_a_type;
  assign T_2006 = io_inner_acquire_bits_is_builtin_type & T_2003;
  assign T_2007 = T_1734 & T_2006;
  assign T_2010 = T_2007 & T_1769;
  assign T_2019 = T_2010 ? 8'hfe : 8'h0;
  assign T_2020 = T_1991 | T_2019;
  assign GEN_32 = T_1962 ? T_2020 : T_175;
  assign GEN_439 = {{3'd0}, 1'h0};
  assign T_2028 = 4'h8 * GEN_439;
  assign T_2030 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_2031 = io_inner_acquire_bits_is_builtin_type & T_2030;
  assign T_2033 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_2034 = io_inner_acquire_bits_is_builtin_type & T_2033;
  assign T_2035 = T_2031 | T_2034;
  assign T_2036 = io_inner_acquire_bits_union[5:1];
  assign T_2037 = T_2035 ? 5'h1 : T_2036;
  assign T_2038 = io_inner_acquire_bits_union[11:9];
  assign T_2039 = io_inner_acquire_bits_union[8:6];
  assign T_2052_0 = 3'h2;
  assign T_2052_1 = 3'h3;
  assign T_2052_2 = 3'h4;
  assign T_2054 = T_2052_0 == io_inner_acquire_bits_a_type;
  assign T_2055 = T_2052_1 == io_inner_acquire_bits_a_type;
  assign T_2056 = T_2052_2 == io_inner_acquire_bits_a_type;
  assign T_2059 = T_2054 | T_2055;
  assign T_2060 = T_2059 | T_2056;
  assign T_2061 = io_inner_acquire_bits_is_builtin_type & T_2060;
  assign T_2062 = T_1734 & T_2061;
  assign GEN_440 = {{7'd0}, T_2062};
  assign T_2064 = 8'h0 - GEN_440;
  assign T_2065 = T_2064[7:0];
  assign T_2066 = ~ T_2065;
  assign T_2070 = T_2066 | T_1989;
  assign T_2072 = T_2034 ? T_2070 : {{7'd0}, 1'h0};
  assign GEN_33 = T_1885 ? io_inner_acquire_bits_addr_block : T_57;
  assign GEN_34 = T_1885 ? 1'h0 : T_59;
  assign GEN_35 = T_1885 ? T_2028 : T_61;
  assign GEN_36 = T_1885 ? T_2037 : T_63;
  assign GEN_37 = T_1885 ? T_2038 : T_65;
  assign GEN_38 = T_1885 ? T_2039 : T_67;
  assign GEN_42 = T_1885 ? T_2072 : GEN_32;
  assign GEN_43 = T_1885 ? {{7'd0}, 1'h0} : T_177;
  assign GEN_44 = T_1885 ? 4'h5 : T_55;
  assign T_2075 = T_175 != GEN_432;
  assign T_2088_0 = 3'h3;
  assign T_2090 = T_2088_0 == T_99_a_type;
  assign T_2093 = T_99_is_builtin_type & T_2090;
  assign T_2094 = T_1887 & T_2093;
  assign T_2095 = T_2094 & T_153;
  assign T_2098 = T_2095 & T_1905;
  assign T_2099 = T_1733 | T_2098;
  assign T_2100 = ~ T_177;
  assign skip_outer_acquire = T_2100 == GEN_432;
  assign T_2109 = 3'h4 == T_99_a_type;
  assign T_2110 = T_2109 ? 2'h0 : 2'h2;
  assign T_2111 = 3'h6 == T_99_a_type;
  assign T_2112 = T_2111 ? 2'h0 : T_2110;
  assign T_2113 = 3'h5 == T_99_a_type;
  assign T_2114 = T_2113 ? 2'h2 : T_2112;
  assign T_2115 = 3'h2 == T_99_a_type;
  assign T_2116 = T_2115 ? 2'h0 : T_2114;
  assign T_2117 = 3'h0 == T_99_a_type;
  assign T_2118 = T_2117 ? 2'h2 : T_2116;
  assign T_2119 = 3'h3 == T_99_a_type;
  assign T_2120 = T_2119 ? 2'h0 : T_2118;
  assign T_2121 = 3'h1 == T_99_a_type;
  assign T_2122 = T_2121 ? 2'h2 : T_2120;
  assign GEN_444 = {{2'd0}, 1'h1};
  assign T_2123 = GEN_444 == T_99_a_type;
  assign T_2124 = T_2123 ? 2'h0 : 2'h2;
  assign T_2125 = GEN_433 == T_99_a_type;
  assign T_2126 = T_2125 ? 2'h1 : T_2124;
  assign T_2127 = T_99_is_builtin_type ? T_2122 : T_2126;
  assign T_2155_addr_block = T_57;
  assign T_2155_p_type = T_2127;
  assign T_2155_client_id = 1'h0;
  assign T_2183 = skip_outer_acquire == 1'h0;
  assign T_2184 = T_2183 ? 4'h6 : 4'h7;
  assign T_2193_pending = T_2276;
  assign T_2193_up_idx = 3'h0;
  assign T_2193_up_done = T_2201;
  assign T_2193_down_idx = T_2259;
  assign T_2193_down_done = T_2260;
  assign T_2201 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2202 = ~ T_2201;
  assign GEN_446 = {{1'd0}, 1'h1};
  assign T_2204 = GEN_446 << io_inner_probe_bits_client_id;
  assign T_2205 = ~ T_2204;
  assign GEN_447 = {{1'd0}, T_2202};
  assign T_2206 = GEN_447 | T_2205;
  assign GEN_448 = {{1'd0}, T_195};
  assign T_2207 = GEN_448 & T_2206;
  assign T_2208 = T_55 == 4'h5;
  assign T_2211 = T_2208 & T_195;
  assign T_2228 = io_inner_release_ready & io_inner_release_valid;
  assign T_2231 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2232 = T_1779 & T_2231;
  assign T_2233 = T_2228 & T_2232;
  assign T_2240_0 = 3'h0;
  assign T_2240_1 = 3'h1;
  assign T_2240_2 = 3'h2;
  assign T_2242 = T_2240_0 == io_inner_release_bits_r_type;
  assign T_2243 = T_2240_1 == io_inner_release_bits_r_type;
  assign T_2244 = T_2240_2 == io_inner_release_bits_r_type;
  assign T_2247 = T_2242 | T_2243;
  assign T_2248 = T_2247 | T_2244;
  assign T_2250 = T_2233 & T_2248;
  assign T_2254 = T_2252 == 3'h7;
  assign T_2256 = T_2252 + GEN_444;
  assign T_2257 = T_2256[2:0];
  assign GEN_46 = T_2250 ? T_2257 : T_2252;
  assign T_2258 = T_2250 & T_2254;
  assign T_2259 = T_2248 ? T_2252 : {{2'd0}, 1'h0};
  assign T_2260 = T_2248 ? T_2258 : T_2233;
  assign T_2264 = T_2260 == 1'h0;
  assign T_2265 = T_2201 & T_2264;
  assign T_2267 = T_2262 + 1'h1;
  assign T_2268 = T_2267[0:0];
  assign GEN_47 = T_2265 ? T_2268 : T_2262;
  assign T_2270 = T_2201 == 1'h0;
  assign T_2271 = T_2260 & T_2270;
  assign T_2273 = T_2262 - 1'h1;
  assign T_2274 = T_2273[0:0];
  assign GEN_48 = T_2271 ? T_2274 : GEN_47;
  assign T_2276 = T_2262 > 1'h0;
  assign T_2280 = T_195 | T_2193_pending;
  assign T_2282 = T_2280 == 1'h0;
  assign T_2283 = T_2208 & T_2282;
  assign GEN_49 = T_2283 ? T_2184 : GEN_44;
  assign T_2287 = T_1733 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2288 = T_2287 & io_inner_release_bits_voluntary;
  assign T_2293 = T_2228 & T_2288;
  assign T_2300_0 = 3'h0;
  assign T_2300_1 = 3'h1;
  assign T_2300_2 = 3'h2;
  assign T_2302 = T_2300_0 == io_inner_release_bits_r_type;
  assign T_2303 = T_2300_1 == io_inner_release_bits_r_type;
  assign T_2304 = T_2300_2 == io_inner_release_bits_r_type;
  assign T_2307 = T_2302 | T_2303;
  assign T_2308 = T_2307 | T_2304;
  assign T_2310 = T_2293 & T_2308;
  assign T_2314 = T_2312 == 3'h7;
  assign T_2316 = T_2312 + GEN_444;
  assign T_2317 = T_2316[2:0];
  assign GEN_50 = T_2310 ? T_2317 : T_2312;
  assign T_2318 = T_2310 & T_2314;
  assign T_2319 = T_2308 ? T_2312 : {{2'd0}, 1'h0};
  assign T_2320 = T_2308 ? T_2318 : T_2293;
  assign T_2321 = io_inner_grant_ready & io_inner_grant_valid;
  assign GEN_452 = {{1'd0}, 3'h0};
  assign T_2324 = io_inner_grant_bits_g_type == GEN_452;
  assign T_2325 = io_inner_grant_bits_is_builtin_type & T_2324;
  assign T_2326 = T_1779 & T_2325;
  assign T_2327 = T_2321 & T_2326;
  assign T_2335_0 = 3'h5;
  assign GEN_453 = {{1'd0}, T_2335_0};
  assign T_2337 = GEN_453 == io_inner_grant_bits_g_type;
  assign T_2345_0 = 2'h0;
  assign T_2345_1 = 2'h1;
  assign GEN_454 = {{2'd0}, T_2345_0};
  assign T_2347 = GEN_454 == io_inner_grant_bits_g_type;
  assign GEN_455 = {{2'd0}, T_2345_1};
  assign T_2348 = GEN_455 == io_inner_grant_bits_g_type;
  assign T_2351 = T_2347 | T_2348;
  assign T_2352 = io_inner_grant_bits_is_builtin_type ? T_2337 : T_2351;
  assign T_2354 = T_2327 & T_2352;
  assign T_2358 = T_2356 == 3'h7;
  assign T_2360 = T_2356 + GEN_444;
  assign T_2361 = T_2360[2:0];
  assign GEN_51 = T_2354 ? T_2361 : T_2356;
  assign T_2362 = T_2354 & T_2358;
  assign T_2363 = T_2352 ? T_2356 : {{2'd0}, 1'h0};
  assign T_2364 = T_2352 ? T_2362 : T_2327;
  assign T_2368 = T_2364 == 1'h0;
  assign T_2369 = T_2320 & T_2368;
  assign T_2371 = T_2366 + 1'h1;
  assign T_2372 = T_2371[0:0];
  assign GEN_52 = T_2369 ? T_2372 : T_2366;
  assign T_2374 = T_2320 == 1'h0;
  assign T_2375 = T_2364 & T_2374;
  assign T_2377 = T_2366 - 1'h1;
  assign T_2378 = T_2377[0:0];
  assign GEN_53 = T_2375 ? T_2378 : GEN_52;
  assign T_2380 = T_2366 > 1'h0;
  assign T_2382 = T_1733 & io_alloc_irel_should;
  assign T_2383 = T_2382 & io_inner_release_valid;
  assign GEN_54 = T_2383 ? io_inner_release_bits_addr_block : GEN_33;
  assign GEN_55 = T_2383 ? 4'h7 : GEN_49;
  assign T_2386 = T_1844 & io_inner_release_bits_voluntary;
  assign T_2392_0 = 4'h0;
  assign T_2392_1 = 4'h8;
  assign T_2394 = T_2392_0 == T_55;
  assign T_2395 = T_2392_1 == T_55;
  assign T_2398 = T_2394 | T_2395;
  assign T_2400 = T_2398 == 1'h0;
  assign T_2401 = T_2386 & T_2400;
  assign T_2403 = T_44 == 1'h0;
  assign T_2404 = T_2401 & T_2403;
  assign T_2405 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2407 = T_2405 == 1'h0;
  assign T_2408 = T_2404 & T_2407;
  assign T_2411 = T_2321 == 1'h0;
  assign T_2412 = T_2408 & T_2411;
  assign T_2414 = T_144_pending == 1'h0;
  assign T_2415 = T_2412 & T_2414;
  assign T_2422_0 = 3'h0;
  assign T_2422_1 = 3'h1;
  assign T_2422_2 = 3'h2;
  assign T_2424 = T_2422_0 == io_inner_release_bits_r_type;
  assign T_2425 = T_2422_1 == io_inner_release_bits_r_type;
  assign T_2426 = T_2422_2 == io_inner_release_bits_r_type;
  assign T_2429 = T_2424 | T_2425;
  assign T_2430 = T_2429 | T_2426;
  assign T_2433 = T_2430 == 1'h0;
  assign T_2435 = io_inner_release_bits_addr_beat == GEN_433;
  assign T_2436 = T_2433 | T_2435;
  assign T_2437 = T_2415 & T_2436;
  assign T_2438 = io_alloc_irel_should | T_2437;
  assign T_2445_0 = 3'h0;
  assign T_2445_1 = 3'h1;
  assign T_2445_2 = 3'h2;
  assign T_2447 = T_2445_0 == io_inner_release_bits_r_type;
  assign T_2448 = T_2445_1 == io_inner_release_bits_r_type;
  assign T_2449 = T_2445_2 == io_inner_release_bits_r_type;
  assign T_2452 = T_2447 | T_2448;
  assign T_2453 = T_2452 | T_2449;
  assign T_2461_0 = 3'h0;
  assign T_2461_1 = 3'h1;
  assign T_2461_2 = 3'h2;
  assign T_2463 = T_2461_0 == io_inner_release_bits_r_type;
  assign T_2464 = T_2461_1 == io_inner_release_bits_r_type;
  assign T_2465 = T_2461_2 == io_inner_release_bits_r_type;
  assign T_2468 = T_2463 | T_2464;
  assign T_2469 = T_2468 | T_2465;
  assign T_2470 = T_2228 & T_2469;
  assign GEN_458 = {{7'd0}, T_2470};
  assign T_2472 = 8'h0 - GEN_458;
  assign T_2473 = T_2472[7:0];
  assign T_2474 = ~ T_2473;
  assign T_2476 = GEN_437 << io_inner_release_bits_addr_beat;
  assign T_2477 = ~ T_2476;
  assign T_2478 = T_2474 | T_2477;
  assign T_2480 = T_2453 ? T_2478 : {{7'd0}, 1'h0};
  assign GEN_56 = T_2438 ? io_inner_release_bits_r_type : T_129;
  assign GEN_57 = T_2438 ? io_inner_release_bits_client_id : T_131;
  assign GEN_58 = T_2438 ? io_inner_release_bits_client_xact_id : T_133;
  assign GEN_65 = T_2438 ? T_2480 : T_135;
  assign T_2484 = T_1844 & T_2231;
  assign T_2486 = T_2484 & T_2208;
  assign T_2488 = T_2438 == 1'h0;
  assign T_2489 = T_2488 & T_2486;
  assign T_2496_0 = 3'h0;
  assign T_2496_1 = 3'h1;
  assign T_2496_2 = 3'h2;
  assign T_2498 = T_2496_0 == io_inner_release_bits_r_type;
  assign T_2499 = T_2496_1 == io_inner_release_bits_r_type;
  assign T_2500 = T_2496_2 == io_inner_release_bits_r_type;
  assign T_2503 = T_2498 | T_2499;
  assign T_2504 = T_2503 | T_2500;
  assign T_2505 = T_2228 & T_2504;
  assign GEN_460 = {{7'd0}, T_2505};
  assign T_2507 = 8'h0 - GEN_460;
  assign T_2508 = T_2507[7:0];
  assign T_2509 = ~ T_2508;
  assign T_2513 = T_2509 | T_2477;
  assign T_2514 = T_135 & T_2513;
  assign GEN_69 = T_2489 ? T_2514 : GEN_65;
  assign GEN_75 = T_2228 ? GEN_56 : T_129;
  assign GEN_76 = T_2228 ? GEN_57 : T_131;
  assign GEN_77 = T_2228 ? GEN_58 : T_133;
  assign GEN_84 = T_2228 ? GEN_69 : T_135;
  assign T_2520_0 = 4'h3;
  assign T_2520_1 = 4'h4;
  assign T_2520_2 = 4'h5;
  assign T_2520_3 = 4'h7;
  assign T_2522 = T_2520_0 == T_55;
  assign T_2523 = T_2520_1 == T_55;
  assign T_2524 = T_2520_2 == T_55;
  assign T_2525 = T_2520_3 == T_55;
  assign T_2528 = T_2522 | T_2523;
  assign T_2529 = T_2528 | T_2524;
  assign T_2530 = T_2529 | T_2525;
  assign T_2531 = T_2530 & T_144_pending;
  assign T_2533 = T_135 != GEN_432;
  assign T_2534 = T_2533 | T_210_pending;
  assign T_2536 = T_2534 == 1'h0;
  assign T_2537 = T_2531 & T_2536;
  assign T_2572_addr_beat = {{2'd0}, 1'h0};
  assign T_2572_addr_block = T_57;
  assign T_2572_client_xact_id = T_133;
  assign T_2572_voluntary = 1'h1;
  assign T_2572_r_type = T_129;
  assign T_2572_data = {{63'd0}, 1'h0};
  assign T_2572_client_id = T_131;
  assign T_2639_addr_beat = {{2'd0}, 1'h0};
  assign T_2639_client_xact_id = T_2572_client_xact_id;
  assign T_2639_manager_xact_id = {{2'd0}, 1'h0};
  assign T_2639_is_builtin_type = 1'h1;
  assign T_2639_g_type = {{1'd0}, 3'h0};
  assign T_2639_data = {{63'd0}, 1'h0};
  assign T_2639_client_id = T_2572_client_id;
  assign T_2679_0 = 4'h0;
  assign T_2679_1 = 4'h8;
  assign T_2681 = T_2679_0 == T_55;
  assign T_2682 = T_2679_1 == T_55;
  assign T_2685 = T_2681 | T_2682;
  assign T_2687 = T_2685 == 1'h0;
  assign T_2688 = T_2386 & T_2687;
  assign T_2691 = T_2688 & T_2403;
  assign T_2695 = T_2691 & T_2407;
  assign T_2699 = T_2695 & T_2411;
  assign T_2702 = T_2699 & T_2414;
  assign T_2709 = T_2702 | T_2486;
  assign T_2716_0 = 3'h0;
  assign T_2716_1 = 3'h1;
  assign T_2716_2 = 3'h2;
  assign T_2718 = T_2716_0 == io_inner_release_bits_r_type;
  assign T_2719 = T_2716_1 == io_inner_release_bits_r_type;
  assign T_2720 = T_2716_2 == io_inner_release_bits_r_type;
  assign T_2723 = T_2718 | T_2719;
  assign T_2724 = T_2723 | T_2720;
  assign T_2725 = T_2228 & T_2724;
  assign GEN_0 = GEN_94;
  assign GEN_88 = GEN_444 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_465 = {{1'd0}, 2'h2};
  assign GEN_89 = GEN_465 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_88;
  assign GEN_466 = {{1'd0}, 2'h3};
  assign GEN_90 = GEN_466 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_89;
  assign GEN_91 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_90;
  assign GEN_92 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_91;
  assign GEN_93 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_92;
  assign GEN_94 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_93;
  assign T_2726 = GEN_0[0];
  assign GEN_1 = GEN_94;
  assign T_2727 = GEN_1[1];
  assign GEN_2 = GEN_94;
  assign T_2728 = GEN_2[2];
  assign GEN_3 = GEN_94;
  assign T_2729 = GEN_3[3];
  assign GEN_4 = GEN_94;
  assign T_2730 = GEN_4[4];
  assign GEN_5 = GEN_94;
  assign T_2731 = GEN_5[5];
  assign GEN_6 = GEN_94;
  assign T_2732 = GEN_6[6];
  assign GEN_7 = GEN_94;
  assign T_2733 = GEN_7[7];
  assign GEN_488 = {{7'd0}, T_2726};
  assign T_2735 = 8'h0 - GEN_488;
  assign T_2736 = T_2735[7:0];
  assign GEN_489 = {{7'd0}, T_2727};
  assign T_2738 = 8'h0 - GEN_489;
  assign T_2739 = T_2738[7:0];
  assign GEN_490 = {{7'd0}, T_2728};
  assign T_2741 = 8'h0 - GEN_490;
  assign T_2742 = T_2741[7:0];
  assign GEN_491 = {{7'd0}, T_2729};
  assign T_2744 = 8'h0 - GEN_491;
  assign T_2745 = T_2744[7:0];
  assign GEN_492 = {{7'd0}, T_2730};
  assign T_2747 = 8'h0 - GEN_492;
  assign T_2748 = T_2747[7:0];
  assign GEN_493 = {{7'd0}, T_2731};
  assign T_2750 = 8'h0 - GEN_493;
  assign T_2751 = T_2750[7:0];
  assign GEN_494 = {{7'd0}, T_2732};
  assign T_2753 = 8'h0 - GEN_494;
  assign T_2754 = T_2753[7:0];
  assign GEN_495 = {{7'd0}, T_2733};
  assign T_2756 = 8'h0 - GEN_495;
  assign T_2757 = T_2756[7:0];
  assign T_2763_0 = T_2736;
  assign T_2763_1 = T_2739;
  assign T_2763_2 = T_2742;
  assign T_2763_3 = T_2745;
  assign T_2763_4 = T_2748;
  assign T_2763_5 = T_2751;
  assign T_2763_6 = T_2754;
  assign T_2763_7 = T_2757;
  assign T_2765 = {T_2763_1,T_2763_0};
  assign T_2766 = {T_2763_3,T_2763_2};
  assign T_2767 = {T_2766,T_2765};
  assign T_2768 = {T_2763_5,T_2763_4};
  assign T_2769 = {T_2763_7,T_2763_6};
  assign T_2770 = {T_2769,T_2768};
  assign T_2771 = {T_2770,T_2767};
  assign T_2772 = ~ T_2771;
  assign T_2773 = T_2772 & io_inner_release_bits_data;
  assign GEN_8 = GEN_150;
  assign GEN_144 = GEN_444 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_145 = GEN_465 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_144;
  assign GEN_146 = GEN_466 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_145;
  assign GEN_147 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_146;
  assign GEN_148 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_147;
  assign GEN_149 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_148;
  assign GEN_150 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_149;
  assign T_2774 = T_2771 & GEN_8;
  assign T_2775 = T_2773 | T_2774;
  assign GEN_9 = T_2775;
  assign GEN_151 = GEN_433 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_152 = GEN_444 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_153 = GEN_465 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_154 = GEN_466 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_155 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_156 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_157 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_158 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_177 = T_2725 ? GEN_151 : data_buffer_0;
  assign GEN_178 = T_2725 ? GEN_152 : data_buffer_1;
  assign GEN_179 = T_2725 ? GEN_153 : data_buffer_2;
  assign GEN_180 = T_2725 ? GEN_154 : data_buffer_3;
  assign GEN_181 = T_2725 ? GEN_155 : data_buffer_4;
  assign GEN_182 = T_2725 ? GEN_156 : data_buffer_5;
  assign GEN_183 = T_2725 ? GEN_157 : data_buffer_6;
  assign GEN_184 = T_2725 ? GEN_158 : data_buffer_7;
  assign T_2806_state = 2'h2;
  assign T_2832 = T_1779 | io_alloc_irel_should;
  assign T_2833 = io_outer_release_ready & io_outer_release_valid;
  assign T_2839_0 = 3'h0;
  assign T_2839_1 = 3'h1;
  assign T_2839_2 = 3'h2;
  assign T_2841 = T_2839_0 == io_outer_release_bits_r_type;
  assign T_2842 = T_2839_1 == io_outer_release_bits_r_type;
  assign T_2843 = T_2839_2 == io_outer_release_bits_r_type;
  assign T_2846 = T_2841 | T_2842;
  assign T_2847 = T_2846 | T_2843;
  assign T_2848 = T_2833 & T_2847;
  assign GEN_503 = {{7'd0}, T_2848};
  assign T_2850 = 8'h0 - GEN_503;
  assign T_2851 = T_2850[7:0];
  assign T_2852 = ~ T_2851;
  assign T_2854 = GEN_437 << io_outer_release_bits_addr_beat;
  assign T_2855 = ~ T_2854;
  assign T_2856 = T_2852 | T_2855;
  assign T_2857 = T_201 & T_2856;
  assign T_2865_0 = 3'h0;
  assign T_2865_1 = 3'h1;
  assign T_2865_2 = 3'h2;
  assign T_2867 = T_2865_0 == io_inner_release_bits_r_type;
  assign T_2868 = T_2865_1 == io_inner_release_bits_r_type;
  assign T_2869 = T_2865_2 == io_inner_release_bits_r_type;
  assign T_2872 = T_2867 | T_2868;
  assign T_2873 = T_2872 | T_2869;
  assign T_2874 = T_2228 & T_2873;
  assign GEN_505 = {{7'd0}, T_2874};
  assign T_2877 = 8'h0 - GEN_505;
  assign T_2878 = T_2877[7:0];
  assign T_2881 = T_2878 & T_2476;
  assign T_2882 = T_2857 | T_2881;
  assign T_2883 = T_2882 | GEN_432;
  assign GEN_191 = T_2832 ? T_2883 : T_201;
  assign GEN_193 = T_2833 ? 1'h0 : T_199;
  assign T_2893 = T_2833 & io_outer_release_bits_voluntary;
  assign T_2900_0 = 3'h0;
  assign T_2900_1 = 3'h1;
  assign T_2900_2 = 3'h2;
  assign T_2902 = T_2900_0 == io_outer_release_bits_r_type;
  assign T_2903 = T_2900_1 == io_outer_release_bits_r_type;
  assign T_2904 = T_2900_2 == io_outer_release_bits_r_type;
  assign T_2907 = T_2902 | T_2903;
  assign T_2908 = T_2907 | T_2904;
  assign T_2910 = T_2893 & T_2908;
  assign T_2914 = T_2912 == 3'h7;
  assign T_2916 = T_2912 + GEN_444;
  assign T_2917 = T_2916[2:0];
  assign GEN_194 = T_2910 ? T_2917 : T_2912;
  assign T_2918 = T_2910 & T_2914;
  assign T_2919 = T_2908 ? T_2912 : {{2'd0}, 1'h0};
  assign T_2920 = T_2908 ? T_2918 : T_2893;
  assign T_2923 = io_outer_grant_bits_g_type == GEN_452;
  assign T_2924 = io_outer_grant_bits_is_builtin_type & T_2923;
  assign T_2925 = T_2405 & T_2924;
  assign T_2933_0 = 3'h5;
  assign GEN_510 = {{1'd0}, T_2933_0};
  assign T_2935 = GEN_510 == io_outer_grant_bits_g_type;
  assign T_2943_0 = 1'h0;
  assign GEN_511 = {{3'd0}, T_2943_0};
  assign T_2945 = GEN_511 == io_outer_grant_bits_g_type;
  assign T_2948 = io_outer_grant_bits_is_builtin_type ? T_2935 : T_2945;
  assign T_2950 = T_2925 & T_2948;
  assign T_2954 = T_2952 == 3'h7;
  assign T_2956 = T_2952 + GEN_444;
  assign T_2957 = T_2956[2:0];
  assign GEN_195 = T_2950 ? T_2957 : T_2952;
  assign T_2958 = T_2950 & T_2954;
  assign T_2959 = T_2948 ? T_2952 : {{2'd0}, 1'h0};
  assign T_2960 = T_2948 ? T_2958 : T_2925;
  assign T_2964 = T_2960 == 1'h0;
  assign T_2965 = T_2920 & T_2964;
  assign T_2967 = T_2962 + 1'h1;
  assign T_2968 = T_2967[0:0];
  assign GEN_196 = T_2965 ? T_2968 : T_2962;
  assign T_2970 = T_2920 == 1'h0;
  assign T_2971 = T_2960 & T_2970;
  assign T_2973 = T_2962 - 1'h1;
  assign T_2974 = T_2973[0:0];
  assign GEN_197 = T_2971 ? T_2974 : GEN_196;
  assign T_2976 = T_2962 > 1'h0;
  assign T_2977 = T_55 == 4'h7;
  assign T_2983_0 = 3'h0;
  assign T_2983_1 = 3'h1;
  assign T_2983_2 = 3'h2;
  assign T_2985 = T_2983_0 == io_outer_release_bits_r_type;
  assign T_2986 = T_2983_1 == io_outer_release_bits_r_type;
  assign T_2987 = T_2983_2 == io_outer_release_bits_r_type;
  assign T_2990 = T_2985 | T_2986;
  assign T_2991 = T_2990 | T_2987;
  assign T_2992 = T_201 >> T_210_up_idx;
  assign T_2993 = T_2992[0];
  assign T_2995 = T_2991 ? T_2993 : T_221;
  assign T_2996 = T_2977 & T_2995;
  assign T_3004_0 = 2'h2;
  assign T_3006 = T_3004_0 == T_2806_state;
  assign T_3009 = T_3006 ? 3'h0 : 3'h3;
  assign T_3045_addr_beat = T_210_up_idx;
  assign T_3045_addr_block = T_57;
  assign T_3045_client_xact_id = {{2'd0}, 1'h0};
  assign T_3045_voluntary = 1'h1;
  assign T_3045_r_type = T_3009;
  assign T_3045_data = GEN_10;
  assign GEN_10 = GEN_204;
  assign GEN_198 = GEN_444 == T_210_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_199 = GEN_465 == T_210_up_idx ? data_buffer_2 : GEN_198;
  assign GEN_200 = GEN_466 == T_210_up_idx ? data_buffer_3 : GEN_199;
  assign GEN_201 = 3'h4 == T_210_up_idx ? data_buffer_4 : GEN_200;
  assign GEN_202 = 3'h5 == T_210_up_idx ? data_buffer_5 : GEN_201;
  assign GEN_203 = 3'h6 == T_210_up_idx ? data_buffer_6 : GEN_202;
  assign GEN_204 = 3'h7 == T_210_up_idx ? data_buffer_7 : GEN_203;
  assign T_3074 = T_99_is_builtin_type == 1'h0;
  assign T_3076 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_3087_0 = 3'h3;
  assign T_3089 = T_3087_0 == io_outer_acquire_bits_a_type;
  assign T_3092 = io_outer_acquire_bits_is_builtin_type & T_3089;
  assign T_3093 = T_3076 & T_3092;
  assign T_3097 = T_3095 == 3'h7;
  assign T_3099 = T_3095 + GEN_444;
  assign T_3100 = T_3099[2:0];
  assign GEN_205 = T_3093 ? T_3100 : T_3095;
  assign T_3101 = T_3093 & T_3097;
  assign T_3102 = T_3092 ? T_3095 : T_69;
  assign T_3103 = T_3092 ? T_3101 : T_3076;
  assign T_3109 = T_2924 == 1'h0;
  assign T_3110 = T_2405 & T_3109;
  assign T_3118_0 = 3'h5;
  assign GEN_518 = {{1'd0}, T_3118_0};
  assign T_3120 = GEN_518 == io_outer_grant_bits_g_type;
  assign T_3128_0 = 1'h0;
  assign GEN_519 = {{3'd0}, T_3128_0};
  assign T_3130 = GEN_519 == io_outer_grant_bits_g_type;
  assign T_3133 = io_outer_grant_bits_is_builtin_type ? T_3120 : T_3130;
  assign T_3135 = T_3110 & T_3133;
  assign T_3139 = T_3137 == 3'h7;
  assign T_3141 = T_3137 + GEN_444;
  assign T_3142 = T_3141[2:0];
  assign GEN_206 = T_3135 ? T_3142 : T_3137;
  assign T_3143 = T_3135 & T_3139;
  assign T_3144 = T_3133 ? T_3137 : T_69;
  assign T_3145 = T_3133 ? T_3143 : T_3110;
  assign T_3149 = T_3145 == 1'h0;
  assign T_3150 = T_3103 & T_3149;
  assign T_3152 = T_3147 + 1'h1;
  assign T_3153 = T_3152[0:0];
  assign GEN_207 = T_3150 ? T_3153 : T_3147;
  assign T_3155 = T_3103 == 1'h0;
  assign T_3156 = T_3145 & T_3155;
  assign T_3158 = T_3147 - 1'h1;
  assign T_3159 = T_3158[0:0];
  assign GEN_208 = T_3156 ? T_3159 : GEN_207;
  assign T_3161 = T_3147 > 1'h0;
  assign T_3162 = T_55 == 4'h6;
  assign T_3163 = T_175 >> T_186_up_idx;
  assign T_3164 = T_3163[0];
  assign T_3166 = T_3164 == 1'h0;
  assign T_3168 = T_59 | T_3166;
  assign T_3169 = T_3162 & T_3168;
  assign T_3172 = T_63 == 5'h1;
  assign T_3173 = T_63 == 5'h7;
  assign T_3174 = T_3172 | T_3173;
  assign T_3175 = T_63[3];
  assign T_3176 = T_63 == 5'h4;
  assign T_3177 = T_3175 | T_3176;
  assign T_3178 = T_3174 | T_3177;
  assign T_3179 = T_63 == 5'h3;
  assign T_3180 = T_3178 | T_3179;
  assign T_3181 = T_63 == 5'h6;
  assign T_3182 = T_3180 | T_3181;
  assign T_3185 = {T_63,1'h1};
  assign T_3216_addr_block = T_57;
  assign T_3216_client_xact_id = {{2'd0}, 1'h0};
  assign T_3216_addr_beat = {{2'd0}, 1'h0};
  assign T_3216_is_builtin_type = 1'h0;
  assign T_3216_a_type = {{2'd0}, T_3182};
  assign T_3216_union = {{6'd0}, T_3185};
  assign T_3216_data = {{63'd0}, 1'h0};
  assign GEN_11 = GEN_215;
  assign GEN_209 = GEN_444 == T_186_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_210 = GEN_465 == T_186_up_idx ? wmask_buffer_2 : GEN_209;
  assign GEN_211 = GEN_466 == T_186_up_idx ? wmask_buffer_3 : GEN_210;
  assign GEN_212 = 3'h4 == T_186_up_idx ? wmask_buffer_4 : GEN_211;
  assign GEN_213 = 3'h5 == T_186_up_idx ? wmask_buffer_5 : GEN_212;
  assign GEN_214 = 3'h6 == T_186_up_idx ? wmask_buffer_6 : GEN_213;
  assign GEN_215 = 3'h7 == T_186_up_idx ? wmask_buffer_7 : GEN_214;
  assign T_3281 = {T_63,1'h0};
  assign T_3282 = {T_65,T_67};
  assign T_3283 = {T_3282,T_3281};
  assign T_3285 = {T_67,T_63};
  assign T_3286 = {T_3285,1'h0};
  assign T_3288 = {GEN_11,1'h0};
  assign T_3300 = T_2111 ? 6'h2 : {{5'd0}, 1'h0};
  assign T_3302 = T_2113 ? 6'h0 : T_3300;
  assign T_3304 = T_2109 ? T_3283 : {{6'd0}, T_3302};
  assign T_3306 = T_2119 ? {{3'd0}, T_3288} : T_3304;
  assign T_3308 = T_2115 ? {{3'd0}, T_3288} : T_3306;
  assign T_3310 = T_2121 ? {{3'd0}, T_3286} : T_3308;
  assign T_3312 = T_2117 ? T_3283 : T_3310;
  assign T_3341_addr_block = T_57;
  assign T_3341_client_xact_id = {{2'd0}, 1'h0};
  assign T_3341_addr_beat = T_186_up_idx;
  assign T_3341_is_builtin_type = 1'h1;
  assign T_3341_a_type = T_99_a_type;
  assign T_3341_union = T_3312;
  assign T_3341_data = GEN_12;
  assign GEN_12 = GEN_222;
  assign GEN_216 = GEN_444 == T_186_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_217 = GEN_465 == T_186_up_idx ? data_buffer_2 : GEN_216;
  assign GEN_218 = GEN_466 == T_186_up_idx ? data_buffer_3 : GEN_217;
  assign GEN_219 = 3'h4 == T_186_up_idx ? data_buffer_4 : GEN_218;
  assign GEN_220 = 3'h5 == T_186_up_idx ? data_buffer_5 : GEN_219;
  assign GEN_221 = 3'h6 == T_186_up_idx ? data_buffer_6 : GEN_220;
  assign GEN_222 = 3'h7 == T_186_up_idx ? data_buffer_7 : GEN_221;
  assign T_3369_addr_block = T_3074 ? T_3216_addr_block : T_3341_addr_block;
  assign T_3369_client_xact_id = T_3074 ? T_3216_client_xact_id : T_3341_client_xact_id;
  assign T_3369_addr_beat = T_3074 ? T_3216_addr_beat : T_3341_addr_beat;
  assign T_3369_is_builtin_type = T_3074 ? T_3216_is_builtin_type : T_3341_is_builtin_type;
  assign T_3369_a_type = T_3074 ? T_3216_a_type : T_3341_a_type;
  assign T_3369_union = T_3074 ? T_3216_union : T_3341_union;
  assign T_3369_data = T_3074 ? T_3216_data : T_3341_data;
  assign T_3398 = T_3162 & T_186_up_done;
  assign GEN_223 = T_3398 ? 4'h7 : GEN_55;
  assign T_3408_0 = 3'h5;
  assign T_3408_1 = 3'h4;
  assign GEN_527 = {{1'd0}, T_3408_0};
  assign T_3410 = GEN_527 == io_outer_grant_bits_g_type;
  assign GEN_528 = {{1'd0}, T_3408_1};
  assign T_3411 = GEN_528 == io_outer_grant_bits_g_type;
  assign T_3414 = T_3410 | T_3411;
  assign T_3420_0 = 1'h0;
  assign GEN_529 = {{3'd0}, T_3420_0};
  assign T_3422 = GEN_529 == io_outer_grant_bits_g_type;
  assign T_3425 = io_outer_grant_bits_is_builtin_type ? T_3414 : T_3422;
  assign T_3426 = T_2405 & T_3425;
  assign GEN_13 = GEN_230;
  assign GEN_224 = GEN_444 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_225 = GEN_465 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_224;
  assign GEN_226 = GEN_466 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_225;
  assign GEN_227 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_226;
  assign GEN_228 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_227;
  assign GEN_229 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_228;
  assign GEN_230 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_229;
  assign T_3427 = GEN_13[0];
  assign GEN_14 = GEN_230;
  assign T_3428 = GEN_14[1];
  assign GEN_15 = GEN_230;
  assign T_3429 = GEN_15[2];
  assign GEN_16 = GEN_230;
  assign T_3430 = GEN_16[3];
  assign GEN_17 = GEN_230;
  assign T_3431 = GEN_17[4];
  assign GEN_18 = GEN_230;
  assign T_3432 = GEN_18[5];
  assign GEN_19 = GEN_230;
  assign T_3433 = GEN_19[6];
  assign GEN_20 = GEN_230;
  assign T_3434 = GEN_20[7];
  assign GEN_554 = {{7'd0}, T_3427};
  assign T_3436 = 8'h0 - GEN_554;
  assign T_3437 = T_3436[7:0];
  assign GEN_555 = {{7'd0}, T_3428};
  assign T_3439 = 8'h0 - GEN_555;
  assign T_3440 = T_3439[7:0];
  assign GEN_556 = {{7'd0}, T_3429};
  assign T_3442 = 8'h0 - GEN_556;
  assign T_3443 = T_3442[7:0];
  assign GEN_557 = {{7'd0}, T_3430};
  assign T_3445 = 8'h0 - GEN_557;
  assign T_3446 = T_3445[7:0];
  assign GEN_558 = {{7'd0}, T_3431};
  assign T_3448 = 8'h0 - GEN_558;
  assign T_3449 = T_3448[7:0];
  assign GEN_559 = {{7'd0}, T_3432};
  assign T_3451 = 8'h0 - GEN_559;
  assign T_3452 = T_3451[7:0];
  assign GEN_560 = {{7'd0}, T_3433};
  assign T_3454 = 8'h0 - GEN_560;
  assign T_3455 = T_3454[7:0];
  assign GEN_561 = {{7'd0}, T_3434};
  assign T_3457 = 8'h0 - GEN_561;
  assign T_3458 = T_3457[7:0];
  assign T_3464_0 = T_3437;
  assign T_3464_1 = T_3440;
  assign T_3464_2 = T_3443;
  assign T_3464_3 = T_3446;
  assign T_3464_4 = T_3449;
  assign T_3464_5 = T_3452;
  assign T_3464_6 = T_3455;
  assign T_3464_7 = T_3458;
  assign T_3466 = {T_3464_1,T_3464_0};
  assign T_3467 = {T_3464_3,T_3464_2};
  assign T_3468 = {T_3467,T_3466};
  assign T_3469 = {T_3464_5,T_3464_4};
  assign T_3470 = {T_3464_7,T_3464_6};
  assign T_3471 = {T_3470,T_3469};
  assign T_3472 = {T_3471,T_3468};
  assign T_3473 = ~ T_3472;
  assign T_3474 = T_3473 & io_outer_grant_bits_data;
  assign GEN_21 = GEN_286;
  assign GEN_280 = GEN_444 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_281 = GEN_465 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_280;
  assign GEN_282 = GEN_466 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_281;
  assign GEN_283 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_282;
  assign GEN_284 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_283;
  assign GEN_285 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_284;
  assign GEN_286 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_285;
  assign T_3475 = T_3472 & GEN_21;
  assign T_3476 = T_3474 | T_3475;
  assign GEN_22 = T_3476;
  assign GEN_287 = GEN_433 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_177;
  assign GEN_288 = GEN_444 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_178;
  assign GEN_289 = GEN_465 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_179;
  assign GEN_290 = GEN_466 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_180;
  assign GEN_291 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_181;
  assign GEN_292 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_182;
  assign GEN_293 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_183;
  assign GEN_294 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_184;
  assign GEN_313 = T_3426 ? GEN_287 : GEN_177;
  assign GEN_314 = T_3426 ? GEN_288 : GEN_178;
  assign GEN_315 = T_3426 ? GEN_289 : GEN_179;
  assign GEN_316 = T_3426 ? GEN_290 : GEN_180;
  assign GEN_317 = T_3426 ? GEN_291 : GEN_181;
  assign GEN_318 = T_3426 ? GEN_292 : GEN_182;
  assign GEN_319 = T_3426 ? GEN_293 : GEN_183;
  assign GEN_320 = T_3426 ? GEN_294 : GEN_184;
  assign T_3477 = T_221 | T_186_pending;
  assign T_3478 = T_3477 | T_210_pending;
  assign T_3489 = T_2325 == 1'h0;
  assign T_3491 = T_2321 & T_3489;
  assign T_3499_0 = 3'h5;
  assign GEN_570 = {{1'd0}, T_3499_0};
  assign T_3501 = GEN_570 == io_inner_grant_bits_g_type;
  assign T_3509_0 = 2'h0;
  assign T_3509_1 = 2'h1;
  assign GEN_571 = {{2'd0}, T_3509_0};
  assign T_3511 = GEN_571 == io_inner_grant_bits_g_type;
  assign GEN_572 = {{2'd0}, T_3509_1};
  assign T_3512 = GEN_572 == io_inner_grant_bits_g_type;
  assign T_3515 = T_3511 | T_3512;
  assign T_3516 = io_inner_grant_bits_is_builtin_type ? T_3501 : T_3515;
  assign T_3518 = T_3491 & T_3516;
  assign T_3522 = T_3520 == 3'h7;
  assign T_3524 = T_3520 + GEN_444;
  assign T_3525 = T_3524[2:0];
  assign GEN_321 = T_3518 ? T_3525 : T_3520;
  assign T_3526 = T_3518 & T_3522;
  assign T_3527 = T_3516 ? T_3520 : {{2'd0}, 1'h0};
  assign T_3528 = T_3516 ? T_3526 : T_3491;
  assign T_3529 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3547 = T_3529 == 1'h0;
  assign T_3548 = T_3528 & T_3547;
  assign T_3550 = T_3545 + 1'h1;
  assign T_3551 = T_3550[0:0];
  assign GEN_323 = T_3548 ? T_3551 : T_3545;
  assign T_3553 = T_3528 == 1'h0;
  assign T_3554 = T_3529 & T_3553;
  assign T_3556 = T_3545 - 1'h1;
  assign T_3557 = T_3556[0:0];
  assign GEN_324 = T_3554 ? T_3557 : GEN_323;
  assign T_3559 = T_3545 > 1'h0;
  assign T_3564 = T_1885 == 1'h0;
  assign T_3573_0 = 3'h5;
  assign T_3573_1 = 3'h4;
  assign GEN_575 = {{1'd0}, T_3573_0};
  assign T_3575 = GEN_575 == io_inner_grant_bits_g_type;
  assign GEN_576 = {{1'd0}, T_3573_1};
  assign T_3576 = GEN_576 == io_inner_grant_bits_g_type;
  assign T_3579 = T_3575 | T_3576;
  assign T_3585_0 = 2'h0;
  assign T_3585_1 = 2'h1;
  assign GEN_577 = {{2'd0}, T_3585_0};
  assign T_3587 = GEN_577 == io_inner_grant_bits_g_type;
  assign GEN_578 = {{2'd0}, T_3585_1};
  assign T_3588 = GEN_578 == io_inner_grant_bits_g_type;
  assign T_3591 = T_3587 | T_3588;
  assign T_3592 = io_inner_grant_bits_is_builtin_type ? T_3579 : T_3591;
  assign T_3593 = T_2321 & T_3592;
  assign GEN_579 = {{7'd0}, T_3593};
  assign T_3595 = 8'h0 - GEN_579;
  assign T_3596 = T_3595[7:0];
  assign T_3597 = ~ T_3596;
  assign T_3599 = GEN_437 << io_inner_grant_bits_addr_beat;
  assign T_3600 = ~ T_3599;
  assign T_3601 = T_3597 | T_3600;
  assign T_3602 = T_177 & T_3601;
  assign T_3610_0 = 3'h0;
  assign T_3610_1 = 3'h1;
  assign T_3610_2 = 3'h2;
  assign T_3612 = T_3610_0 == io_inner_release_bits_r_type;
  assign T_3613 = T_3610_1 == io_inner_release_bits_r_type;
  assign T_3614 = T_3610_2 == io_inner_release_bits_r_type;
  assign T_3617 = T_3612 | T_3613;
  assign T_3618 = T_3617 | T_3614;
  assign T_3619 = T_2228 & T_3618;
  assign GEN_581 = {{7'd0}, T_3619};
  assign T_3622 = 8'h0 - GEN_581;
  assign T_3623 = T_3622[7:0];
  assign T_3626 = T_3623 & T_2476;
  assign T_3627 = T_3602 | T_3626;
  assign T_3637_0 = 3'h5;
  assign T_3637_1 = 3'h4;
  assign GEN_583 = {{1'd0}, T_3637_0};
  assign T_3639 = GEN_583 == io_outer_grant_bits_g_type;
  assign GEN_584 = {{1'd0}, T_3637_1};
  assign T_3640 = GEN_584 == io_outer_grant_bits_g_type;
  assign T_3643 = T_3639 | T_3640;
  assign T_3649_0 = 1'h0;
  assign GEN_585 = {{3'd0}, T_3649_0};
  assign T_3651 = GEN_585 == io_outer_grant_bits_g_type;
  assign T_3654 = io_outer_grant_bits_is_builtin_type ? T_3643 : T_3651;
  assign T_3655 = T_2405 & T_3654;
  assign GEN_586 = {{7'd0}, T_3655};
  assign T_3658 = 8'h0 - GEN_586;
  assign T_3659 = T_3658[7:0];
  assign T_3661 = GEN_437 << io_outer_grant_bits_addr_beat;
  assign T_3662 = T_3659 & T_3661;
  assign T_3663 = T_3627 | T_3662;
  assign T_3664 = T_3663 | GEN_432;
  assign GEN_335 = T_3564 ? T_3664 : GEN_43;
  assign T_3666 = T_55 == 4'h1;
  assign T_3667 = T_1733 | T_3666;
  assign T_3670 = T_3667 | T_2075;
  assign T_3672 = T_3670 == 1'h0;
  assign T_3689 = 3'h6 == Queue_11_1_io_deq_bits_a_type;
  assign T_3690 = T_3689 ? 3'h1 : 3'h3;
  assign T_3691 = 3'h5 == Queue_11_1_io_deq_bits_a_type;
  assign T_3692 = T_3691 ? 3'h1 : T_3690;
  assign T_3693 = 3'h4 == Queue_11_1_io_deq_bits_a_type;
  assign T_3694 = T_3693 ? 3'h4 : T_3692;
  assign T_3695 = 3'h3 == Queue_11_1_io_deq_bits_a_type;
  assign T_3696 = T_3695 ? 3'h3 : T_3694;
  assign T_3697 = 3'h2 == Queue_11_1_io_deq_bits_a_type;
  assign T_3698 = T_3697 ? 3'h3 : T_3696;
  assign T_3699 = 3'h1 == Queue_11_1_io_deq_bits_a_type;
  assign T_3700 = T_3699 ? 3'h5 : T_3698;
  assign T_3701 = 3'h0 == Queue_11_1_io_deq_bits_a_type;
  assign T_3702 = T_3701 ? 3'h4 : T_3700;
  assign T_3703 = Queue_11_1_io_deq_bits_a_type == GEN_433;
  assign T_3708 = T_3703 ? 2'h0 : 2'h1;
  assign T_3709 = Queue_11_1_io_deq_bits_is_builtin_type ? T_3702 : {{1'd0}, T_3708};
  assign T_3741_addr_beat = Queue_11_1_io_deq_bits_addr_beat;
  assign T_3741_client_xact_id = Queue_11_1_io_deq_bits_client_xact_id;
  assign T_3741_manager_xact_id = {{2'd0}, 1'h1};
  assign T_3741_is_builtin_type = Queue_11_1_io_deq_bits_is_builtin_type;
  assign T_3741_g_type = {{1'd0}, T_3709};
  assign T_3741_data = GEN_23;
  assign T_3741_client_id = Queue_11_1_io_deq_bits_client_id;
  assign GEN_23 = GEN_342;
  assign GEN_336 = GEN_444 == T_155 ? data_buffer_1 : data_buffer_0;
  assign GEN_337 = GEN_465 == T_155 ? data_buffer_2 : GEN_336;
  assign GEN_338 = GEN_466 == T_155 ? data_buffer_3 : GEN_337;
  assign GEN_339 = 3'h4 == T_155 ? data_buffer_4 : GEN_338;
  assign GEN_340 = 3'h5 == T_155 ? data_buffer_5 : GEN_339;
  assign GEN_341 = 3'h6 == T_155 ? data_buffer_6 : GEN_340;
  assign GEN_342 = 3'h7 == T_155 ? data_buffer_7 : GEN_341;
  assign T_3780_0 = 3'h5;
  assign GEN_594 = {{1'd0}, T_3780_0};
  assign T_3782 = GEN_594 == io_inner_grant_bits_g_type;
  assign T_3790_0 = 2'h0;
  assign T_3790_1 = 2'h1;
  assign GEN_595 = {{2'd0}, T_3790_0};
  assign T_3792 = GEN_595 == io_inner_grant_bits_g_type;
  assign GEN_596 = {{2'd0}, T_3790_1};
  assign T_3793 = GEN_596 == io_inner_grant_bits_g_type;
  assign T_3796 = T_3792 | T_3793;
  assign T_3797 = io_inner_grant_bits_is_builtin_type ? T_3782 : T_3796;
  assign T_3799 = T_2321 & T_3797;
  assign T_3803 = T_3801 == 3'h7;
  assign T_3805 = T_3801 + GEN_444;
  assign T_3806 = T_3805[2:0];
  assign GEN_343 = T_3799 ? T_3806 : T_3801;
  assign T_3807 = T_3799 & T_3803;
  assign T_3808 = T_3797 ? T_3801 : Queue_11_1_io_deq_bits_addr_beat;
  assign T_3809 = T_3797 ? T_3807 : T_2321;
  assign T_3814 = T_2977 & T_153;
  assign T_3816 = T_3478 == 1'h0;
  assign T_3824_0 = 3'h5;
  assign T_3824_1 = 3'h4;
  assign GEN_598 = {{1'd0}, T_3824_0};
  assign T_3826 = GEN_598 == io_inner_grant_bits_g_type;
  assign GEN_599 = {{1'd0}, T_3824_1};
  assign T_3827 = GEN_599 == io_inner_grant_bits_g_type;
  assign T_3830 = T_3826 | T_3827;
  assign T_3836_0 = 2'h0;
  assign T_3836_1 = 2'h1;
  assign GEN_600 = {{2'd0}, T_3836_0};
  assign T_3838 = GEN_600 == io_inner_grant_bits_g_type;
  assign GEN_601 = {{2'd0}, T_3836_1};
  assign T_3839 = GEN_601 == io_inner_grant_bits_g_type;
  assign T_3842 = T_3838 | T_3839;
  assign T_3843 = io_inner_grant_bits_is_builtin_type ? T_3830 : T_3842;
  assign T_3844 = T_177 >> T_155;
  assign T_3845 = T_3844[0];
  assign T_3846 = T_3843 ? T_3845 : T_3672;
  assign T_3847 = T_3816 & T_3846;
  assign GEN_348 = T_3814 ? T_3847 : T_2537;
  assign GEN_349 = T_2414 ? T_157 : 1'h0;
  assign GEN_350 = T_2414 ? T_155 : T_2639_addr_beat;
  assign GEN_351 = T_2414 ? T_3741_client_xact_id : T_2639_client_xact_id;
  assign GEN_352 = T_2414 ? T_3741_manager_xact_id : T_2639_manager_xact_id;
  assign GEN_353 = T_2414 ? T_3741_is_builtin_type : T_2639_is_builtin_type;
  assign GEN_354 = T_2414 ? T_3741_g_type : T_2639_g_type;
  assign GEN_355 = T_2414 ? T_3741_data : T_2639_data;
  assign GEN_356 = T_2414 ? T_3741_client_id : T_2639_client_id;
  assign GEN_361 = T_2414 ? GEN_348 : T_2537;
  assign T_3854 = ~ io_incoherent_0;
  assign GEN_362 = T_1885 ? {{1'd0}, T_3854} : T_2207;
  assign T_3869_0 = 3'h3;
  assign T_3871 = T_3869_0 == T_99_a_type;
  assign T_3874 = T_99_is_builtin_type & T_3871;
  assign T_3875 = T_1887 & T_3874;
  assign T_3876 = T_3875 & T_153;
  assign T_3879 = T_3876 & T_1905;
  assign T_3881 = T_3879 & io_inner_acquire_valid;
  assign T_3882 = T_1885 | T_3881;
  assign T_3892_0 = 3'h2;
  assign T_3892_1 = 3'h3;
  assign T_3892_2 = 3'h4;
  assign T_3894 = T_3892_0 == io_inner_acquire_bits_a_type;
  assign T_3895 = T_3892_1 == io_inner_acquire_bits_a_type;
  assign T_3896 = T_3892_2 == io_inner_acquire_bits_a_type;
  assign T_3899 = T_3894 | T_3895;
  assign T_3900 = T_3899 | T_3896;
  assign T_3901 = io_inner_acquire_bits_is_builtin_type & T_3900;
  assign T_3902 = T_1734 & T_3901;
  assign T_3903 = T_3902 & T_3882;
  assign T_3905 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3906 = io_inner_acquire_bits_is_builtin_type & T_3905;
  assign T_3910 = 8'h0 - GEN_437;
  assign T_3911 = T_3910[7:0];
  assign T_3917_0 = T_3911;
  assign T_3925 = T_2034 | T_2031;
  assign T_3926 = io_inner_acquire_bits_union[8:1];
  assign T_3928 = T_3925 ? T_3926 : {{7'd0}, 1'h0};
  assign T_3929 = T_3906 ? T_3917_0 : T_3928;
  assign T_3930 = T_3929[0];
  assign T_3931 = T_3929[1];
  assign T_3932 = T_3929[2];
  assign T_3933 = T_3929[3];
  assign T_3934 = T_3929[4];
  assign T_3935 = T_3929[5];
  assign T_3936 = T_3929[6];
  assign T_3937 = T_3929[7];
  assign GEN_603 = {{7'd0}, T_3930};
  assign T_3939 = 8'h0 - GEN_603;
  assign T_3940 = T_3939[7:0];
  assign GEN_604 = {{7'd0}, T_3931};
  assign T_3942 = 8'h0 - GEN_604;
  assign T_3943 = T_3942[7:0];
  assign GEN_605 = {{7'd0}, T_3932};
  assign T_3945 = 8'h0 - GEN_605;
  assign T_3946 = T_3945[7:0];
  assign GEN_606 = {{7'd0}, T_3933};
  assign T_3948 = 8'h0 - GEN_606;
  assign T_3949 = T_3948[7:0];
  assign GEN_607 = {{7'd0}, T_3934};
  assign T_3951 = 8'h0 - GEN_607;
  assign T_3952 = T_3951[7:0];
  assign GEN_608 = {{7'd0}, T_3935};
  assign T_3954 = 8'h0 - GEN_608;
  assign T_3955 = T_3954[7:0];
  assign GEN_609 = {{7'd0}, T_3936};
  assign T_3957 = 8'h0 - GEN_609;
  assign T_3958 = T_3957[7:0];
  assign GEN_610 = {{7'd0}, T_3937};
  assign T_3960 = 8'h0 - GEN_610;
  assign T_3961 = T_3960[7:0];
  assign T_3967_0 = T_3940;
  assign T_3967_1 = T_3943;
  assign T_3967_2 = T_3946;
  assign T_3967_3 = T_3949;
  assign T_3967_4 = T_3952;
  assign T_3967_5 = T_3955;
  assign T_3967_6 = T_3958;
  assign T_3967_7 = T_3961;
  assign T_3969 = {T_3967_1,T_3967_0};
  assign T_3970 = {T_3967_3,T_3967_2};
  assign T_3971 = {T_3970,T_3969};
  assign T_3972 = {T_3967_5,T_3967_4};
  assign T_3973 = {T_3967_7,T_3967_6};
  assign T_3974 = {T_3973,T_3972};
  assign T_3975 = {T_3974,T_3971};
  assign T_3976 = ~ T_3975;
  assign GEN_24 = GEN_369;
  assign GEN_363 = GEN_444 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_364 = GEN_465 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_363;
  assign GEN_365 = GEN_466 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_364;
  assign GEN_366 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_365;
  assign GEN_367 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_366;
  assign GEN_368 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_367;
  assign GEN_369 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_368;
  assign T_3977 = T_3976 & GEN_24;
  assign T_3978 = T_3975 & io_inner_acquire_bits_data;
  assign T_3979 = T_3977 | T_3978;
  assign GEN_25 = T_3979;
  assign GEN_370 = GEN_433 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_313;
  assign GEN_371 = GEN_444 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_314;
  assign GEN_372 = GEN_465 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_315;
  assign GEN_373 = GEN_466 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_316;
  assign GEN_374 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_317;
  assign GEN_375 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_318;
  assign GEN_376 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_319;
  assign GEN_377 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_320;
  assign T_3993_0 = T_3911;
  assign T_4005 = T_3906 ? T_3993_0 : T_3928;
  assign GEN_26 = GEN_384;
  assign GEN_378 = GEN_444 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_379 = GEN_465 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_378;
  assign GEN_380 = GEN_466 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_379;
  assign GEN_381 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_380;
  assign GEN_382 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_381;
  assign GEN_383 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_382;
  assign GEN_384 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_383;
  assign T_4006 = T_4005 | GEN_26;
  assign GEN_27 = T_4006;
  assign GEN_385 = GEN_433 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_0;
  assign GEN_386 = GEN_444 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_1;
  assign GEN_387 = GEN_465 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_2;
  assign GEN_388 = GEN_466 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_3;
  assign GEN_389 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_4;
  assign GEN_390 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_5;
  assign GEN_391 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_6;
  assign GEN_392 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_7;
  assign GEN_404 = T_3903 ? GEN_370 : GEN_313;
  assign GEN_405 = T_3903 ? GEN_371 : GEN_314;
  assign GEN_406 = T_3903 ? GEN_372 : GEN_315;
  assign GEN_407 = T_3903 ? GEN_373 : GEN_316;
  assign GEN_408 = T_3903 ? GEN_374 : GEN_317;
  assign GEN_409 = T_3903 ? GEN_375 : GEN_318;
  assign GEN_410 = T_3903 ? GEN_376 : GEN_319;
  assign GEN_411 = T_3903 ? GEN_377 : GEN_320;
  assign GEN_415 = T_3903 ? GEN_385 : wmask_buffer_0;
  assign GEN_416 = T_3903 ? GEN_386 : wmask_buffer_1;
  assign GEN_417 = T_3903 ? GEN_387 : wmask_buffer_2;
  assign GEN_418 = T_3903 ? GEN_388 : wmask_buffer_3;
  assign GEN_419 = T_3903 ? GEN_389 : wmask_buffer_4;
  assign GEN_420 = T_3903 ? GEN_390 : wmask_buffer_5;
  assign GEN_421 = T_3903 ? GEN_391 : wmask_buffer_6;
  assign GEN_422 = T_3903 ? GEN_392 : wmask_buffer_7;
  assign T_4009 = T_2075 | T_2533;
  assign T_4010 = T_4009 | T_144_pending;
  assign T_4011 = T_4010 | T_221;
  assign T_4012 = T_4011 | T_210_pending;
  assign T_4013 = T_4012 | T_186_pending;
  assign T_4014 = T_4013 | T_153;
  assign T_4015 = T_4014 | T_166_pending;
  assign T_4017 = T_4015 == 1'h0;
  assign T_4019 = T_2977 & T_44;
  assign GEN_423 = T_4019 ? 4'h0 : GEN_223;
  assign GEN_424 = T_4019 ? {{7'd0}, 1'h0} : GEN_415;
  assign GEN_425 = T_4019 ? {{7'd0}, 1'h0} : GEN_416;
  assign GEN_426 = T_4019 ? {{7'd0}, 1'h0} : GEN_417;
  assign GEN_427 = T_4019 ? {{7'd0}, 1'h0} : GEN_418;
  assign GEN_428 = T_4019 ? {{7'd0}, 1'h0} : GEN_419;
  assign GEN_429 = T_4019 ? {{7'd0}, 1'h0} : GEN_420;
  assign GEN_430 = T_4019 ? {{7'd0}, 1'h0} : GEN_421;
  assign GEN_431 = T_4019 ? {{7'd0}, 1'h0} : GEN_422;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_30 = {1{$random}};
  T_55 = GEN_30[3:0];
  GEN_31 = {1{$random}};
  T_57 = GEN_31[25:0];
  GEN_39 = {1{$random}};
  T_59 = GEN_39[0:0];
  GEN_40 = {1{$random}};
  T_61 = GEN_40[4:0];
  GEN_41 = {1{$random}};
  T_63 = GEN_41[4:0];
  GEN_45 = {1{$random}};
  T_65 = GEN_45[2:0];
  GEN_59 = {1{$random}};
  T_67 = GEN_59[2:0];
  GEN_60 = {1{$random}};
  T_129 = GEN_60[2:0];
  GEN_61 = {1{$random}};
  T_131 = GEN_61[0:0];
  GEN_62 = {1{$random}};
  T_133 = GEN_62[1:0];
  GEN_63 = {1{$random}};
  T_135 = GEN_63[7:0];
  GEN_64 = {1{$random}};
  T_175 = GEN_64[7:0];
  GEN_66 = {1{$random}};
  T_177 = GEN_66[7:0];
  GEN_67 = {1{$random}};
  T_195 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  T_199 = GEN_68[0:0];
  GEN_70 = {1{$random}};
  T_201 = GEN_70[7:0];
  GEN_71 = {2{$random}};
  data_buffer_0 = GEN_71[63:0];
  GEN_72 = {2{$random}};
  data_buffer_1 = GEN_72[63:0];
  GEN_73 = {2{$random}};
  data_buffer_2 = GEN_73[63:0];
  GEN_74 = {2{$random}};
  data_buffer_3 = GEN_74[63:0];
  GEN_78 = {2{$random}};
  data_buffer_4 = GEN_78[63:0];
  GEN_79 = {2{$random}};
  data_buffer_5 = GEN_79[63:0];
  GEN_80 = {2{$random}};
  data_buffer_6 = GEN_80[63:0];
  GEN_81 = {2{$random}};
  data_buffer_7 = GEN_81[63:0];
  GEN_82 = {1{$random}};
  wmask_buffer_0 = GEN_82[7:0];
  GEN_83 = {1{$random}};
  wmask_buffer_1 = GEN_83[7:0];
  GEN_85 = {1{$random}};
  wmask_buffer_2 = GEN_85[7:0];
  GEN_86 = {1{$random}};
  wmask_buffer_3 = GEN_86[7:0];
  GEN_87 = {1{$random}};
  wmask_buffer_4 = GEN_87[7:0];
  GEN_95 = {1{$random}};
  wmask_buffer_5 = GEN_95[7:0];
  GEN_96 = {1{$random}};
  wmask_buffer_6 = GEN_96[7:0];
  GEN_97 = {1{$random}};
  wmask_buffer_7 = GEN_97[7:0];
  GEN_98 = {1{$random}};
  T_2219 = GEN_98[2:0];
  GEN_99 = {1{$random}};
  T_2252 = GEN_99[2:0];
  GEN_100 = {1{$random}};
  T_2262 = GEN_100[0:0];
  GEN_101 = {1{$random}};
  T_2312 = GEN_101[2:0];
  GEN_102 = {1{$random}};
  T_2356 = GEN_102[2:0];
  GEN_103 = {1{$random}};
  T_2366 = GEN_103[0:0];
  GEN_104 = {1{$random}};
  T_2912 = GEN_104[2:0];
  GEN_105 = {1{$random}};
  T_2952 = GEN_105[2:0];
  GEN_106 = {1{$random}};
  T_2962 = GEN_106[0:0];
  GEN_107 = {1{$random}};
  T_3095 = GEN_107[2:0];
  GEN_108 = {1{$random}};
  T_3137 = GEN_108[2:0];
  GEN_109 = {1{$random}};
  T_3147 = GEN_109[0:0];
  GEN_110 = {1{$random}};
  T_3520 = GEN_110[2:0];
  GEN_111 = {1{$random}};
  T_3535 = GEN_111[2:0];
  GEN_112 = {1{$random}};
  T_3545 = GEN_112[0:0];
  GEN_113 = {1{$random}};
  T_3801 = GEN_113[2:0];
  GEN_114 = {1{$random}};
  GEN_28 = GEN_114[0:0];
  GEN_115 = {1{$random}};
  GEN_29 = GEN_115[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_55 <= 4'h0;
    end else begin
      if(T_4019) begin
        T_55 <= 4'h0;
      end else begin
        if(T_3398) begin
          T_55 <= 4'h7;
        end else begin
          if(T_2383) begin
            T_55 <= 4'h7;
          end else begin
            if(T_2283) begin
              if(T_2183) begin
                T_55 <= 4'h6;
              end else begin
                T_55 <= 4'h7;
              end
            end else begin
              if(T_1885) begin
                T_55 <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_57 <= 26'h0;
    end else begin
      if(T_2383) begin
        T_57 <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1885) begin
          T_57 <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_59 <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_61 <= T_2028;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        if(T_2035) begin
          T_63 <= 5'h1;
        end else begin
          T_63 <= T_2036;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_65 <= T_2038;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_67 <= T_2039;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_129 <= io_inner_release_bits_r_type;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_131 <= io_inner_release_bits_client_id;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_133 <= io_inner_release_bits_client_xact_id;
        end
      end
    end
    if(reset) begin
      T_135 <= 8'h0;
    end else begin
      if(T_2228) begin
        if(T_2489) begin
          T_135 <= T_2514;
        end else begin
          if(T_2438) begin
            if(T_2453) begin
              T_135 <= T_2478;
            end else begin
              T_135 <= {{7'd0}, 1'h0};
            end
          end
        end
      end
    end
    if(reset) begin
      T_175 <= 8'h0;
    end else begin
      if(T_1885) begin
        if(T_2034) begin
          T_175 <= T_2070;
        end else begin
          T_175 <= {{7'd0}, 1'h0};
        end
      end else begin
        if(T_1962) begin
          T_175 <= T_2020;
        end
      end
    end
    if(reset) begin
      T_177 <= 8'h0;
    end else begin
      if(T_3564) begin
        T_177 <= T_3664;
      end else begin
        if(T_1885) begin
          T_177 <= {{7'd0}, 1'h0};
        end
      end
    end
    if(1'h0) begin
    end else begin
      T_195 <= GEN_362[0];
    end
    if(reset) begin
      T_199 <= 1'h0;
    end else begin
      if(T_2833) begin
        T_199 <= 1'h0;
      end
    end
    if(reset) begin
      T_201 <= 8'h0;
    end else begin
      if(T_2832) begin
        T_201 <= T_2883;
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1817_0;
    end else begin
      if(T_3903) begin
        if(GEN_433 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_433 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_433 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_433 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_433 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_433 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_433 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1817_1;
    end else begin
      if(T_3903) begin
        if(GEN_444 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_444 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_444 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_444 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_444 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_444 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_444 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1817_2;
    end else begin
      if(T_3903) begin
        if(GEN_465 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_465 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_465 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_465 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_465 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_465 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_465 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1817_3;
    end else begin
      if(T_3903) begin
        if(GEN_466 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_466 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_466 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_466 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_466 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_466 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_466 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1817_4;
    end else begin
      if(T_3903) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1817_5;
    end else begin
      if(T_3903) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1817_6;
    end else begin
      if(T_3903) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1817_7;
    end else begin
      if(T_3903) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1835_0;
    end else begin
      if(T_4019) begin
        wmask_buffer_0 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_433 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1835_1;
    end else begin
      if(T_4019) begin
        wmask_buffer_1 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_444 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1835_2;
    end else begin
      if(T_4019) begin
        wmask_buffer_2 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_465 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1835_3;
    end else begin
      if(T_4019) begin
        wmask_buffer_3 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_466 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1835_4;
    end else begin
      if(T_4019) begin
        wmask_buffer_4 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1835_5;
    end else begin
      if(T_4019) begin
        wmask_buffer_5 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1835_6;
    end else begin
      if(T_4019) begin
        wmask_buffer_6 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1835_7;
    end else begin
      if(T_4019) begin
        wmask_buffer_7 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      T_2219 <= 3'h0;
    end
    if(reset) begin
      T_2252 <= 3'h0;
    end else begin
      if(T_2250) begin
        T_2252 <= T_2257;
      end
    end
    if(reset) begin
      T_2262 <= 1'h0;
    end else begin
      if(T_2271) begin
        T_2262 <= T_2274;
      end else begin
        if(T_2265) begin
          T_2262 <= T_2268;
        end
      end
    end
    if(reset) begin
      T_2312 <= 3'h0;
    end else begin
      if(T_2310) begin
        T_2312 <= T_2317;
      end
    end
    if(reset) begin
      T_2356 <= 3'h0;
    end else begin
      if(T_2354) begin
        T_2356 <= T_2361;
      end
    end
    if(reset) begin
      T_2366 <= 1'h0;
    end else begin
      if(T_2375) begin
        T_2366 <= T_2378;
      end else begin
        if(T_2369) begin
          T_2366 <= T_2372;
        end
      end
    end
    if(reset) begin
      T_2912 <= 3'h0;
    end else begin
      if(T_2910) begin
        T_2912 <= T_2917;
      end
    end
    if(reset) begin
      T_2952 <= 3'h0;
    end else begin
      if(T_2950) begin
        T_2952 <= T_2957;
      end
    end
    if(reset) begin
      T_2962 <= 1'h0;
    end else begin
      if(T_2971) begin
        T_2962 <= T_2974;
      end else begin
        if(T_2965) begin
          T_2962 <= T_2968;
        end
      end
    end
    if(reset) begin
      T_3095 <= 3'h0;
    end else begin
      if(T_3093) begin
        T_3095 <= T_3100;
      end
    end
    if(reset) begin
      T_3137 <= 3'h0;
    end else begin
      if(T_3135) begin
        T_3137 <= T_3142;
      end
    end
    if(reset) begin
      T_3147 <= 1'h0;
    end else begin
      if(T_3156) begin
        T_3147 <= T_3159;
      end else begin
        if(T_3150) begin
          T_3147 <= T_3153;
        end
      end
    end
    if(reset) begin
      T_3520 <= 3'h0;
    end else begin
      if(T_3518) begin
        T_3520 <= T_3525;
      end
    end
    if(reset) begin
      T_3535 <= 3'h0;
    end
    if(reset) begin
      T_3545 <= 1'h0;
    end else begin
      if(T_3554) begin
        T_3545 <= T_3557;
      end else begin
        if(T_3548) begin
          T_3545 <= T_3551;
        end
      end
    end
    if(reset) begin
      T_3801 <= 3'h0;
    end else begin
      if(T_3799) begin
        T_3801 <= T_3806;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1778) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:95 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1778) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1778) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1792) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:99 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1792) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1792) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1803) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1803) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1803) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BufferedBroadcastAcquireTracker_1(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should
);
  wire  T_44;
  reg [3:0] T_55;
  reg [31:0] GEN_30;
  reg [25:0] T_57;
  reg [31:0] GEN_31;
  reg  T_59;
  reg [31:0] GEN_39;
  reg [4:0] T_61;
  reg [31:0] GEN_40;
  reg [4:0] T_63;
  reg [31:0] GEN_41;
  reg [2:0] T_65;
  reg [31:0] GEN_45;
  reg [2:0] T_67;
  reg [31:0] GEN_59;
  wire [2:0] T_69;
  wire [1:0] T_99_client_xact_id;
  wire [2:0] T_99_addr_beat;
  wire  T_99_client_id;
  wire  T_99_is_builtin_type;
  wire [2:0] T_99_a_type;
  reg [2:0] T_129;
  reg [31:0] GEN_60;
  reg  T_131;
  reg [31:0] GEN_61;
  reg [1:0] T_133;
  reg [31:0] GEN_62;
  reg [7:0] T_135;
  reg [31:0] GEN_63;
  wire  T_144_pending;
  wire [2:0] T_144_up_idx;
  wire  T_144_up_done;
  wire [2:0] T_144_down_idx;
  wire  T_144_down_done;
  wire  T_153;
  wire [2:0] T_155;
  wire  T_157;
  wire  T_166_pending;
  wire [2:0] T_166_up_idx;
  wire  T_166_up_done;
  wire [2:0] T_166_down_idx;
  wire  T_166_down_done;
  reg [7:0] T_175;
  reg [31:0] GEN_64;
  reg [7:0] T_177;
  reg [31:0] GEN_66;
  wire  T_186_pending;
  wire [2:0] T_186_up_idx;
  wire  T_186_up_done;
  wire [2:0] T_186_down_idx;
  wire  T_186_down_done;
  reg  T_195;
  reg [31:0] GEN_67;
  reg  T_199;
  reg [31:0] GEN_68;
  reg [7:0] T_201;
  reg [31:0] GEN_70;
  wire  T_210_pending;
  wire [2:0] T_210_up_idx;
  wire  T_210_up_done;
  wire [2:0] T_210_down_idx;
  wire  T_210_down_done;
  wire [7:0] GEN_432;
  wire  T_219;
  wire  T_220;
  wire  T_221;
  wire  T_247_sharers;
  wire [1:0] T_299_state;
  wire  T_395_inner_sharers;
  wire [1:0] T_395_outer_state;
  wire  T_1733;
  wire  T_1734;
  wire  T_1735;
  wire  T_1736;
  wire [2:0] T_1745_0;
  wire  T_1747;
  wire  T_1750;
  wire  T_1751;
  wire [2:0] T_1760_0;
  wire  T_1762;
  wire  T_1765;
  wire  T_1767;
  wire [2:0] GEN_433;
  wire  T_1769;
  wire  T_1770;
  wire  T_1772;
  wire  T_1773;
  wire  T_1775;
  wire  T_1776;
  wire  T_1778;
  wire  T_1779;
  wire  T_1780;
  wire  T_1782;
  wire  T_1784;
  wire  T_1785;
  wire  T_1786;
  wire  T_1787;
  wire  T_1789;
  wire  T_1790;
  wire  T_1792;
  wire  T_1796;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [63:0] T_1817_0;
  wire [63:0] T_1817_1;
  wire [63:0] T_1817_2;
  wire [63:0] T_1817_3;
  wire [63:0] T_1817_4;
  wire [63:0] T_1817_5;
  wire [63:0] T_1817_6;
  wire [63:0] T_1817_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_71;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_72;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_73;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_74;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_78;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_79;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_80;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_81;
  wire [7:0] T_1835_0;
  wire [7:0] T_1835_1;
  wire [7:0] T_1835_2;
  wire [7:0] T_1835_3;
  wire [7:0] T_1835_4;
  wire [7:0] T_1835_5;
  wire [7:0] T_1835_6;
  wire [7:0] T_1835_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_82;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_83;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_85;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_86;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_87;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_95;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_96;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_97;
  wire  T_1841;
  wire  T_1842;
  wire  T_1844;
  wire  T_1845;
  wire  T_1847;
  wire  T_1848;
  wire  Queue_12_1_clk;
  wire  Queue_12_1_reset;
  wire  Queue_12_1_io_enq_ready;
  wire  Queue_12_1_io_enq_valid;
  wire [1:0] Queue_12_1_io_enq_bits_client_xact_id;
  wire [2:0] Queue_12_1_io_enq_bits_addr_beat;
  wire  Queue_12_1_io_enq_bits_client_id;
  wire  Queue_12_1_io_enq_bits_is_builtin_type;
  wire [2:0] Queue_12_1_io_enq_bits_a_type;
  wire  Queue_12_1_io_deq_ready;
  wire  Queue_12_1_io_deq_valid;
  wire [1:0] Queue_12_1_io_deq_bits_client_xact_id;
  wire [2:0] Queue_12_1_io_deq_bits_addr_beat;
  wire  Queue_12_1_io_deq_bits_client_id;
  wire  Queue_12_1_io_deq_bits_is_builtin_type;
  wire [2:0] Queue_12_1_io_deq_bits_a_type;
  wire [1:0] Queue_12_1_io_count;
  wire  T_1884;
  wire  T_1885;
  wire  T_1887;
  wire [2:0] T_1896_0;
  wire  T_1898;
  wire  T_1901;
  wire  T_1902;
  wire  T_1903;
  wire [7:0] T_1904;
  wire  T_1905;
  wire  T_1906;
  wire  T_1908;
  wire [2:0] T_1917_0;
  wire  T_1919;
  wire  T_1922;
  wire  T_1924;
  wire  T_1927;
  wire  T_1928;
  wire  T_1929;
  wire [1:0] T_1930_client_xact_id;
  wire [2:0] T_1930_addr_beat;
  wire  T_1930_client_id;
  wire  T_1930_is_builtin_type;
  wire [2:0] T_1930_a_type;
  wire [1:0] GEN_435;
  wire  T_1960;
  wire  T_1962;
  wire [2:0] T_1972_0;
  wire [2:0] T_1972_1;
  wire [2:0] T_1972_2;
  wire  T_1974;
  wire  T_1975;
  wire  T_1976;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire  T_1982;
  wire [7:0] GEN_436;
  wire [8:0] T_1984;
  wire [7:0] T_1985;
  wire [7:0] T_1986;
  wire [7:0] GEN_437;
  wire [7:0] T_1988;
  wire [7:0] T_1989;
  wire [7:0] T_1990;
  wire [7:0] T_1991;
  wire [2:0] T_2001_0;
  wire  T_2003;
  wire  T_2006;
  wire  T_2007;
  wire  T_2010;
  wire [7:0] T_2019;
  wire [7:0] T_2020;
  wire [7:0] GEN_32;
  wire [3:0] GEN_439;
  wire [4:0] T_2028;
  wire  T_2030;
  wire  T_2031;
  wire  T_2033;
  wire  T_2034;
  wire  T_2035;
  wire [4:0] T_2036;
  wire [4:0] T_2037;
  wire [2:0] T_2038;
  wire [2:0] T_2039;
  wire [2:0] T_2052_0;
  wire [2:0] T_2052_1;
  wire [2:0] T_2052_2;
  wire  T_2054;
  wire  T_2055;
  wire  T_2056;
  wire  T_2059;
  wire  T_2060;
  wire  T_2061;
  wire  T_2062;
  wire [7:0] GEN_440;
  wire [8:0] T_2064;
  wire [7:0] T_2065;
  wire [7:0] T_2066;
  wire [7:0] T_2070;
  wire [7:0] T_2072;
  wire [25:0] GEN_33;
  wire  GEN_34;
  wire [4:0] GEN_35;
  wire [4:0] GEN_36;
  wire [2:0] GEN_37;
  wire [2:0] GEN_38;
  wire [7:0] GEN_42;
  wire [7:0] GEN_43;
  wire [3:0] GEN_44;
  wire  T_2075;
  wire [2:0] T_2088_0;
  wire  T_2090;
  wire  T_2093;
  wire  T_2094;
  wire  T_2095;
  wire  T_2098;
  wire  T_2099;
  wire [7:0] T_2100;
  wire  skip_outer_acquire;
  wire  T_2109;
  wire [1:0] T_2110;
  wire  T_2111;
  wire [1:0] T_2112;
  wire  T_2113;
  wire [1:0] T_2114;
  wire  T_2115;
  wire [1:0] T_2116;
  wire  T_2117;
  wire [1:0] T_2118;
  wire  T_2119;
  wire [1:0] T_2120;
  wire  T_2121;
  wire [1:0] T_2122;
  wire [2:0] GEN_444;
  wire  T_2123;
  wire [1:0] T_2124;
  wire  T_2125;
  wire [1:0] T_2126;
  wire [1:0] T_2127;
  wire [25:0] T_2155_addr_block;
  wire [1:0] T_2155_p_type;
  wire  T_2155_client_id;
  wire  T_2183;
  wire [3:0] T_2184;
  wire  T_2193_pending;
  wire [2:0] T_2193_up_idx;
  wire  T_2193_up_done;
  wire [2:0] T_2193_down_idx;
  wire  T_2193_down_done;
  wire  T_2201;
  wire  T_2202;
  wire [1:0] GEN_446;
  wire [1:0] T_2204;
  wire [1:0] T_2205;
  wire [1:0] GEN_447;
  wire [1:0] T_2206;
  wire [1:0] GEN_448;
  wire [1:0] T_2207;
  wire  T_2208;
  wire  T_2211;
  reg [2:0] T_2219;
  reg [31:0] GEN_98;
  wire  T_2228;
  wire  T_2231;
  wire  T_2232;
  wire  T_2233;
  wire [2:0] T_2240_0;
  wire [2:0] T_2240_1;
  wire [2:0] T_2240_2;
  wire  T_2242;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  reg [2:0] T_2252;
  reg [31:0] GEN_99;
  wire  T_2254;
  wire [3:0] T_2256;
  wire [2:0] T_2257;
  wire [2:0] GEN_46;
  wire  T_2258;
  wire [2:0] T_2259;
  wire  T_2260;
  reg  T_2262;
  reg [31:0] GEN_100;
  wire  T_2264;
  wire  T_2265;
  wire [1:0] T_2267;
  wire  T_2268;
  wire  GEN_47;
  wire  T_2270;
  wire  T_2271;
  wire [1:0] T_2273;
  wire  T_2274;
  wire  GEN_48;
  wire  T_2276;
  wire  T_2280;
  wire  T_2282;
  wire  T_2283;
  wire [3:0] GEN_49;
  wire  T_2287;
  wire  T_2288;
  wire  T_2293;
  wire [2:0] T_2300_0;
  wire [2:0] T_2300_1;
  wire [2:0] T_2300_2;
  wire  T_2302;
  wire  T_2303;
  wire  T_2304;
  wire  T_2307;
  wire  T_2308;
  wire  T_2310;
  reg [2:0] T_2312;
  reg [31:0] GEN_101;
  wire  T_2314;
  wire [3:0] T_2316;
  wire [2:0] T_2317;
  wire [2:0] GEN_50;
  wire  T_2318;
  wire [2:0] T_2319;
  wire  T_2320;
  wire  T_2321;
  wire [3:0] GEN_452;
  wire  T_2324;
  wire  T_2325;
  wire  T_2326;
  wire  T_2327;
  wire [2:0] T_2335_0;
  wire [3:0] GEN_453;
  wire  T_2337;
  wire [1:0] T_2345_0;
  wire [1:0] T_2345_1;
  wire [3:0] GEN_454;
  wire  T_2347;
  wire [3:0] GEN_455;
  wire  T_2348;
  wire  T_2351;
  wire  T_2352;
  wire  T_2354;
  reg [2:0] T_2356;
  reg [31:0] GEN_102;
  wire  T_2358;
  wire [3:0] T_2360;
  wire [2:0] T_2361;
  wire [2:0] GEN_51;
  wire  T_2362;
  wire [2:0] T_2363;
  wire  T_2364;
  reg  T_2366;
  reg [31:0] GEN_103;
  wire  T_2368;
  wire  T_2369;
  wire [1:0] T_2371;
  wire  T_2372;
  wire  GEN_52;
  wire  T_2374;
  wire  T_2375;
  wire [1:0] T_2377;
  wire  T_2378;
  wire  GEN_53;
  wire  T_2380;
  wire  T_2382;
  wire  T_2383;
  wire [25:0] GEN_54;
  wire [3:0] GEN_55;
  wire  T_2386;
  wire [3:0] T_2392_0;
  wire [3:0] T_2392_1;
  wire  T_2394;
  wire  T_2395;
  wire  T_2398;
  wire  T_2400;
  wire  T_2401;
  wire  T_2403;
  wire  T_2404;
  wire  T_2405;
  wire  T_2407;
  wire  T_2408;
  wire  T_2411;
  wire  T_2412;
  wire  T_2414;
  wire  T_2415;
  wire [2:0] T_2422_0;
  wire [2:0] T_2422_1;
  wire [2:0] T_2422_2;
  wire  T_2424;
  wire  T_2425;
  wire  T_2426;
  wire  T_2429;
  wire  T_2430;
  wire  T_2433;
  wire  T_2435;
  wire  T_2436;
  wire  T_2437;
  wire  T_2438;
  wire [2:0] T_2445_0;
  wire [2:0] T_2445_1;
  wire [2:0] T_2445_2;
  wire  T_2447;
  wire  T_2448;
  wire  T_2449;
  wire  T_2452;
  wire  T_2453;
  wire [2:0] T_2461_0;
  wire [2:0] T_2461_1;
  wire [2:0] T_2461_2;
  wire  T_2463;
  wire  T_2464;
  wire  T_2465;
  wire  T_2468;
  wire  T_2469;
  wire  T_2470;
  wire [7:0] GEN_458;
  wire [8:0] T_2472;
  wire [7:0] T_2473;
  wire [7:0] T_2474;
  wire [7:0] T_2476;
  wire [7:0] T_2477;
  wire [7:0] T_2478;
  wire [7:0] T_2480;
  wire [2:0] GEN_56;
  wire  GEN_57;
  wire [1:0] GEN_58;
  wire [7:0] GEN_65;
  wire  T_2484;
  wire  T_2486;
  wire  T_2488;
  wire  T_2489;
  wire [2:0] T_2496_0;
  wire [2:0] T_2496_1;
  wire [2:0] T_2496_2;
  wire  T_2498;
  wire  T_2499;
  wire  T_2500;
  wire  T_2503;
  wire  T_2504;
  wire  T_2505;
  wire [7:0] GEN_460;
  wire [8:0] T_2507;
  wire [7:0] T_2508;
  wire [7:0] T_2509;
  wire [7:0] T_2513;
  wire [7:0] T_2514;
  wire [7:0] GEN_69;
  wire [2:0] GEN_75;
  wire  GEN_76;
  wire [1:0] GEN_77;
  wire [7:0] GEN_84;
  wire [3:0] T_2520_0;
  wire [3:0] T_2520_1;
  wire [3:0] T_2520_2;
  wire [3:0] T_2520_3;
  wire  T_2522;
  wire  T_2523;
  wire  T_2524;
  wire  T_2525;
  wire  T_2528;
  wire  T_2529;
  wire  T_2530;
  wire  T_2531;
  wire  T_2533;
  wire  T_2534;
  wire  T_2536;
  wire  T_2537;
  wire [2:0] T_2572_addr_beat;
  wire [25:0] T_2572_addr_block;
  wire [1:0] T_2572_client_xact_id;
  wire  T_2572_voluntary;
  wire [2:0] T_2572_r_type;
  wire [63:0] T_2572_data;
  wire  T_2572_client_id;
  wire [2:0] T_2639_addr_beat;
  wire [1:0] T_2639_client_xact_id;
  wire [2:0] T_2639_manager_xact_id;
  wire  T_2639_is_builtin_type;
  wire [3:0] T_2639_g_type;
  wire [63:0] T_2639_data;
  wire  T_2639_client_id;
  wire [3:0] T_2679_0;
  wire [3:0] T_2679_1;
  wire  T_2681;
  wire  T_2682;
  wire  T_2685;
  wire  T_2687;
  wire  T_2688;
  wire  T_2691;
  wire  T_2695;
  wire  T_2699;
  wire  T_2702;
  wire  T_2709;
  wire [2:0] T_2716_0;
  wire [2:0] T_2716_1;
  wire [2:0] T_2716_2;
  wire  T_2718;
  wire  T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [7:0] GEN_0;
  wire [7:0] GEN_88;
  wire [2:0] GEN_465;
  wire [7:0] GEN_89;
  wire [2:0] GEN_466;
  wire [7:0] GEN_90;
  wire [7:0] GEN_91;
  wire [7:0] GEN_92;
  wire [7:0] GEN_93;
  wire [7:0] GEN_94;
  wire  T_2726;
  wire [7:0] GEN_1;
  wire  T_2727;
  wire [7:0] GEN_2;
  wire  T_2728;
  wire [7:0] GEN_3;
  wire  T_2729;
  wire [7:0] GEN_4;
  wire  T_2730;
  wire [7:0] GEN_5;
  wire  T_2731;
  wire [7:0] GEN_6;
  wire  T_2732;
  wire [7:0] GEN_7;
  wire  T_2733;
  wire [7:0] GEN_488;
  wire [8:0] T_2735;
  wire [7:0] T_2736;
  wire [7:0] GEN_489;
  wire [8:0] T_2738;
  wire [7:0] T_2739;
  wire [7:0] GEN_490;
  wire [8:0] T_2741;
  wire [7:0] T_2742;
  wire [7:0] GEN_491;
  wire [8:0] T_2744;
  wire [7:0] T_2745;
  wire [7:0] GEN_492;
  wire [8:0] T_2747;
  wire [7:0] T_2748;
  wire [7:0] GEN_493;
  wire [8:0] T_2750;
  wire [7:0] T_2751;
  wire [7:0] GEN_494;
  wire [8:0] T_2753;
  wire [7:0] T_2754;
  wire [7:0] GEN_495;
  wire [8:0] T_2756;
  wire [7:0] T_2757;
  wire [7:0] T_2763_0;
  wire [7:0] T_2763_1;
  wire [7:0] T_2763_2;
  wire [7:0] T_2763_3;
  wire [7:0] T_2763_4;
  wire [7:0] T_2763_5;
  wire [7:0] T_2763_6;
  wire [7:0] T_2763_7;
  wire [15:0] T_2765;
  wire [15:0] T_2766;
  wire [31:0] T_2767;
  wire [15:0] T_2768;
  wire [15:0] T_2769;
  wire [31:0] T_2770;
  wire [63:0] T_2771;
  wire [63:0] T_2772;
  wire [63:0] T_2773;
  wire [63:0] GEN_8;
  wire [63:0] GEN_144;
  wire [63:0] GEN_145;
  wire [63:0] GEN_146;
  wire [63:0] GEN_147;
  wire [63:0] GEN_148;
  wire [63:0] GEN_149;
  wire [63:0] GEN_150;
  wire [63:0] T_2774;
  wire [63:0] T_2775;
  wire [63:0] GEN_9;
  wire [63:0] GEN_151;
  wire [63:0] GEN_152;
  wire [63:0] GEN_153;
  wire [63:0] GEN_154;
  wire [63:0] GEN_155;
  wire [63:0] GEN_156;
  wire [63:0] GEN_157;
  wire [63:0] GEN_158;
  wire [63:0] GEN_177;
  wire [63:0] GEN_178;
  wire [63:0] GEN_179;
  wire [63:0] GEN_180;
  wire [63:0] GEN_181;
  wire [63:0] GEN_182;
  wire [63:0] GEN_183;
  wire [63:0] GEN_184;
  wire [1:0] T_2806_state;
  wire  T_2832;
  wire  T_2833;
  wire [2:0] T_2839_0;
  wire [2:0] T_2839_1;
  wire [2:0] T_2839_2;
  wire  T_2841;
  wire  T_2842;
  wire  T_2843;
  wire  T_2846;
  wire  T_2847;
  wire  T_2848;
  wire [7:0] GEN_503;
  wire [8:0] T_2850;
  wire [7:0] T_2851;
  wire [7:0] T_2852;
  wire [7:0] T_2854;
  wire [7:0] T_2855;
  wire [7:0] T_2856;
  wire [7:0] T_2857;
  wire [2:0] T_2865_0;
  wire [2:0] T_2865_1;
  wire [2:0] T_2865_2;
  wire  T_2867;
  wire  T_2868;
  wire  T_2869;
  wire  T_2872;
  wire  T_2873;
  wire  T_2874;
  wire [7:0] GEN_505;
  wire [8:0] T_2877;
  wire [7:0] T_2878;
  wire [7:0] T_2881;
  wire [7:0] T_2882;
  wire [7:0] T_2883;
  wire [7:0] GEN_191;
  wire  GEN_193;
  wire  T_2893;
  wire [2:0] T_2900_0;
  wire [2:0] T_2900_1;
  wire [2:0] T_2900_2;
  wire  T_2902;
  wire  T_2903;
  wire  T_2904;
  wire  T_2907;
  wire  T_2908;
  wire  T_2910;
  reg [2:0] T_2912;
  reg [31:0] GEN_104;
  wire  T_2914;
  wire [3:0] T_2916;
  wire [2:0] T_2917;
  wire [2:0] GEN_194;
  wire  T_2918;
  wire [2:0] T_2919;
  wire  T_2920;
  wire  T_2923;
  wire  T_2924;
  wire  T_2925;
  wire [2:0] T_2933_0;
  wire [3:0] GEN_510;
  wire  T_2935;
  wire  T_2943_0;
  wire [3:0] GEN_511;
  wire  T_2945;
  wire  T_2948;
  wire  T_2950;
  reg [2:0] T_2952;
  reg [31:0] GEN_105;
  wire  T_2954;
  wire [3:0] T_2956;
  wire [2:0] T_2957;
  wire [2:0] GEN_195;
  wire  T_2958;
  wire [2:0] T_2959;
  wire  T_2960;
  reg  T_2962;
  reg [31:0] GEN_106;
  wire  T_2964;
  wire  T_2965;
  wire [1:0] T_2967;
  wire  T_2968;
  wire  GEN_196;
  wire  T_2970;
  wire  T_2971;
  wire [1:0] T_2973;
  wire  T_2974;
  wire  GEN_197;
  wire  T_2976;
  wire  T_2977;
  wire [2:0] T_2983_0;
  wire [2:0] T_2983_1;
  wire [2:0] T_2983_2;
  wire  T_2985;
  wire  T_2986;
  wire  T_2987;
  wire  T_2990;
  wire  T_2991;
  wire [7:0] T_2992;
  wire  T_2993;
  wire  T_2995;
  wire  T_2996;
  wire [1:0] T_3004_0;
  wire  T_3006;
  wire [2:0] T_3009;
  wire [2:0] T_3045_addr_beat;
  wire [25:0] T_3045_addr_block;
  wire [2:0] T_3045_client_xact_id;
  wire  T_3045_voluntary;
  wire [2:0] T_3045_r_type;
  wire [63:0] T_3045_data;
  wire [63:0] GEN_10;
  wire [63:0] GEN_198;
  wire [63:0] GEN_199;
  wire [63:0] GEN_200;
  wire [63:0] GEN_201;
  wire [63:0] GEN_202;
  wire [63:0] GEN_203;
  wire [63:0] GEN_204;
  wire  T_3074;
  wire  T_3076;
  wire [2:0] T_3087_0;
  wire  T_3089;
  wire  T_3092;
  wire  T_3093;
  reg [2:0] T_3095;
  reg [31:0] GEN_107;
  wire  T_3097;
  wire [3:0] T_3099;
  wire [2:0] T_3100;
  wire [2:0] GEN_205;
  wire  T_3101;
  wire [2:0] T_3102;
  wire  T_3103;
  wire  T_3109;
  wire  T_3110;
  wire [2:0] T_3118_0;
  wire [3:0] GEN_518;
  wire  T_3120;
  wire  T_3128_0;
  wire [3:0] GEN_519;
  wire  T_3130;
  wire  T_3133;
  wire  T_3135;
  reg [2:0] T_3137;
  reg [31:0] GEN_108;
  wire  T_3139;
  wire [3:0] T_3141;
  wire [2:0] T_3142;
  wire [2:0] GEN_206;
  wire  T_3143;
  wire [2:0] T_3144;
  wire  T_3145;
  reg  T_3147;
  reg [31:0] GEN_109;
  wire  T_3149;
  wire  T_3150;
  wire [1:0] T_3152;
  wire  T_3153;
  wire  GEN_207;
  wire  T_3155;
  wire  T_3156;
  wire [1:0] T_3158;
  wire  T_3159;
  wire  GEN_208;
  wire  T_3161;
  wire  T_3162;
  wire [7:0] T_3163;
  wire  T_3164;
  wire  T_3166;
  wire  T_3168;
  wire  T_3169;
  wire  T_3172;
  wire  T_3173;
  wire  T_3174;
  wire  T_3175;
  wire  T_3176;
  wire  T_3177;
  wire  T_3178;
  wire  T_3179;
  wire  T_3180;
  wire  T_3181;
  wire  T_3182;
  wire [5:0] T_3185;
  wire [25:0] T_3216_addr_block;
  wire [2:0] T_3216_client_xact_id;
  wire [2:0] T_3216_addr_beat;
  wire  T_3216_is_builtin_type;
  wire [2:0] T_3216_a_type;
  wire [11:0] T_3216_union;
  wire [63:0] T_3216_data;
  wire [7:0] GEN_11;
  wire [7:0] GEN_209;
  wire [7:0] GEN_210;
  wire [7:0] GEN_211;
  wire [7:0] GEN_212;
  wire [7:0] GEN_213;
  wire [7:0] GEN_214;
  wire [7:0] GEN_215;
  wire [5:0] T_3281;
  wire [5:0] T_3282;
  wire [11:0] T_3283;
  wire [7:0] T_3285;
  wire [8:0] T_3286;
  wire [8:0] T_3288;
  wire [5:0] T_3300;
  wire [5:0] T_3302;
  wire [11:0] T_3304;
  wire [11:0] T_3306;
  wire [11:0] T_3308;
  wire [11:0] T_3310;
  wire [11:0] T_3312;
  wire [25:0] T_3341_addr_block;
  wire [2:0] T_3341_client_xact_id;
  wire [2:0] T_3341_addr_beat;
  wire  T_3341_is_builtin_type;
  wire [2:0] T_3341_a_type;
  wire [11:0] T_3341_union;
  wire [63:0] T_3341_data;
  wire [63:0] GEN_12;
  wire [63:0] GEN_216;
  wire [63:0] GEN_217;
  wire [63:0] GEN_218;
  wire [63:0] GEN_219;
  wire [63:0] GEN_220;
  wire [63:0] GEN_221;
  wire [63:0] GEN_222;
  wire [25:0] T_3369_addr_block;
  wire [2:0] T_3369_client_xact_id;
  wire [2:0] T_3369_addr_beat;
  wire  T_3369_is_builtin_type;
  wire [2:0] T_3369_a_type;
  wire [11:0] T_3369_union;
  wire [63:0] T_3369_data;
  wire  T_3398;
  wire [3:0] GEN_223;
  wire [2:0] T_3408_0;
  wire [2:0] T_3408_1;
  wire [3:0] GEN_527;
  wire  T_3410;
  wire [3:0] GEN_528;
  wire  T_3411;
  wire  T_3414;
  wire  T_3420_0;
  wire [3:0] GEN_529;
  wire  T_3422;
  wire  T_3425;
  wire  T_3426;
  wire [7:0] GEN_13;
  wire [7:0] GEN_224;
  wire [7:0] GEN_225;
  wire [7:0] GEN_226;
  wire [7:0] GEN_227;
  wire [7:0] GEN_228;
  wire [7:0] GEN_229;
  wire [7:0] GEN_230;
  wire  T_3427;
  wire [7:0] GEN_14;
  wire  T_3428;
  wire [7:0] GEN_15;
  wire  T_3429;
  wire [7:0] GEN_16;
  wire  T_3430;
  wire [7:0] GEN_17;
  wire  T_3431;
  wire [7:0] GEN_18;
  wire  T_3432;
  wire [7:0] GEN_19;
  wire  T_3433;
  wire [7:0] GEN_20;
  wire  T_3434;
  wire [7:0] GEN_554;
  wire [8:0] T_3436;
  wire [7:0] T_3437;
  wire [7:0] GEN_555;
  wire [8:0] T_3439;
  wire [7:0] T_3440;
  wire [7:0] GEN_556;
  wire [8:0] T_3442;
  wire [7:0] T_3443;
  wire [7:0] GEN_557;
  wire [8:0] T_3445;
  wire [7:0] T_3446;
  wire [7:0] GEN_558;
  wire [8:0] T_3448;
  wire [7:0] T_3449;
  wire [7:0] GEN_559;
  wire [8:0] T_3451;
  wire [7:0] T_3452;
  wire [7:0] GEN_560;
  wire [8:0] T_3454;
  wire [7:0] T_3455;
  wire [7:0] GEN_561;
  wire [8:0] T_3457;
  wire [7:0] T_3458;
  wire [7:0] T_3464_0;
  wire [7:0] T_3464_1;
  wire [7:0] T_3464_2;
  wire [7:0] T_3464_3;
  wire [7:0] T_3464_4;
  wire [7:0] T_3464_5;
  wire [7:0] T_3464_6;
  wire [7:0] T_3464_7;
  wire [15:0] T_3466;
  wire [15:0] T_3467;
  wire [31:0] T_3468;
  wire [15:0] T_3469;
  wire [15:0] T_3470;
  wire [31:0] T_3471;
  wire [63:0] T_3472;
  wire [63:0] T_3473;
  wire [63:0] T_3474;
  wire [63:0] GEN_21;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [63:0] GEN_286;
  wire [63:0] T_3475;
  wire [63:0] T_3476;
  wire [63:0] GEN_22;
  wire [63:0] GEN_287;
  wire [63:0] GEN_288;
  wire [63:0] GEN_289;
  wire [63:0] GEN_290;
  wire [63:0] GEN_291;
  wire [63:0] GEN_292;
  wire [63:0] GEN_293;
  wire [63:0] GEN_294;
  wire [63:0] GEN_313;
  wire [63:0] GEN_314;
  wire [63:0] GEN_315;
  wire [63:0] GEN_316;
  wire [63:0] GEN_317;
  wire [63:0] GEN_318;
  wire [63:0] GEN_319;
  wire [63:0] GEN_320;
  wire  T_3477;
  wire  T_3478;
  wire  T_3489;
  wire  T_3491;
  wire [2:0] T_3499_0;
  wire [3:0] GEN_570;
  wire  T_3501;
  wire [1:0] T_3509_0;
  wire [1:0] T_3509_1;
  wire [3:0] GEN_571;
  wire  T_3511;
  wire [3:0] GEN_572;
  wire  T_3512;
  wire  T_3515;
  wire  T_3516;
  wire  T_3518;
  reg [2:0] T_3520;
  reg [31:0] GEN_110;
  wire  T_3522;
  wire [3:0] T_3524;
  wire [2:0] T_3525;
  wire [2:0] GEN_321;
  wire  T_3526;
  wire [2:0] T_3527;
  wire  T_3528;
  wire  T_3529;
  reg [2:0] T_3535;
  reg [31:0] GEN_111;
  reg  T_3545;
  reg [31:0] GEN_112;
  wire  T_3547;
  wire  T_3548;
  wire [1:0] T_3550;
  wire  T_3551;
  wire  GEN_323;
  wire  T_3553;
  wire  T_3554;
  wire [1:0] T_3556;
  wire  T_3557;
  wire  GEN_324;
  wire  T_3559;
  wire  T_3564;
  wire [2:0] T_3573_0;
  wire [2:0] T_3573_1;
  wire [3:0] GEN_575;
  wire  T_3575;
  wire [3:0] GEN_576;
  wire  T_3576;
  wire  T_3579;
  wire [1:0] T_3585_0;
  wire [1:0] T_3585_1;
  wire [3:0] GEN_577;
  wire  T_3587;
  wire [3:0] GEN_578;
  wire  T_3588;
  wire  T_3591;
  wire  T_3592;
  wire  T_3593;
  wire [7:0] GEN_579;
  wire [8:0] T_3595;
  wire [7:0] T_3596;
  wire [7:0] T_3597;
  wire [7:0] T_3599;
  wire [7:0] T_3600;
  wire [7:0] T_3601;
  wire [7:0] T_3602;
  wire [2:0] T_3610_0;
  wire [2:0] T_3610_1;
  wire [2:0] T_3610_2;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3617;
  wire  T_3618;
  wire  T_3619;
  wire [7:0] GEN_581;
  wire [8:0] T_3622;
  wire [7:0] T_3623;
  wire [7:0] T_3626;
  wire [7:0] T_3627;
  wire [2:0] T_3637_0;
  wire [2:0] T_3637_1;
  wire [3:0] GEN_583;
  wire  T_3639;
  wire [3:0] GEN_584;
  wire  T_3640;
  wire  T_3643;
  wire  T_3649_0;
  wire [3:0] GEN_585;
  wire  T_3651;
  wire  T_3654;
  wire  T_3655;
  wire [7:0] GEN_586;
  wire [8:0] T_3658;
  wire [7:0] T_3659;
  wire [7:0] T_3661;
  wire [7:0] T_3662;
  wire [7:0] T_3663;
  wire [7:0] T_3664;
  wire [7:0] GEN_335;
  wire  T_3666;
  wire  T_3667;
  wire  T_3670;
  wire  T_3672;
  wire  T_3689;
  wire [2:0] T_3690;
  wire  T_3691;
  wire [2:0] T_3692;
  wire  T_3693;
  wire [2:0] T_3694;
  wire  T_3695;
  wire [2:0] T_3696;
  wire  T_3697;
  wire [2:0] T_3698;
  wire  T_3699;
  wire [2:0] T_3700;
  wire  T_3701;
  wire [2:0] T_3702;
  wire  T_3703;
  wire [1:0] T_3708;
  wire [2:0] T_3709;
  wire [2:0] T_3741_addr_beat;
  wire [1:0] T_3741_client_xact_id;
  wire [2:0] T_3741_manager_xact_id;
  wire  T_3741_is_builtin_type;
  wire [3:0] T_3741_g_type;
  wire [63:0] T_3741_data;
  wire  T_3741_client_id;
  wire [63:0] GEN_23;
  wire [63:0] GEN_336;
  wire [63:0] GEN_337;
  wire [63:0] GEN_338;
  wire [63:0] GEN_339;
  wire [63:0] GEN_340;
  wire [63:0] GEN_341;
  wire [63:0] GEN_342;
  wire [2:0] T_3780_0;
  wire [3:0] GEN_594;
  wire  T_3782;
  wire [1:0] T_3790_0;
  wire [1:0] T_3790_1;
  wire [3:0] GEN_595;
  wire  T_3792;
  wire [3:0] GEN_596;
  wire  T_3793;
  wire  T_3796;
  wire  T_3797;
  wire  T_3799;
  reg [2:0] T_3801;
  reg [31:0] GEN_113;
  wire  T_3803;
  wire [3:0] T_3805;
  wire [2:0] T_3806;
  wire [2:0] GEN_343;
  wire  T_3807;
  wire [2:0] T_3808;
  wire  T_3809;
  wire  T_3814;
  wire  T_3816;
  wire [2:0] T_3824_0;
  wire [2:0] T_3824_1;
  wire [3:0] GEN_598;
  wire  T_3826;
  wire [3:0] GEN_599;
  wire  T_3827;
  wire  T_3830;
  wire [1:0] T_3836_0;
  wire [1:0] T_3836_1;
  wire [3:0] GEN_600;
  wire  T_3838;
  wire [3:0] GEN_601;
  wire  T_3839;
  wire  T_3842;
  wire  T_3843;
  wire [7:0] T_3844;
  wire  T_3845;
  wire  T_3846;
  wire  T_3847;
  wire  GEN_348;
  wire  GEN_349;
  wire [2:0] GEN_350;
  wire [1:0] GEN_351;
  wire [2:0] GEN_352;
  wire  GEN_353;
  wire [3:0] GEN_354;
  wire [63:0] GEN_355;
  wire  GEN_356;
  wire  GEN_361;
  wire  T_3854;
  wire [1:0] GEN_362;
  wire [2:0] T_3869_0;
  wire  T_3871;
  wire  T_3874;
  wire  T_3875;
  wire  T_3876;
  wire  T_3879;
  wire  T_3881;
  wire  T_3882;
  wire [2:0] T_3892_0;
  wire [2:0] T_3892_1;
  wire [2:0] T_3892_2;
  wire  T_3894;
  wire  T_3895;
  wire  T_3896;
  wire  T_3899;
  wire  T_3900;
  wire  T_3901;
  wire  T_3902;
  wire  T_3903;
  wire  T_3905;
  wire  T_3906;
  wire [8:0] T_3910;
  wire [7:0] T_3911;
  wire [7:0] T_3917_0;
  wire  T_3925;
  wire [7:0] T_3926;
  wire [7:0] T_3928;
  wire [7:0] T_3929;
  wire  T_3930;
  wire  T_3931;
  wire  T_3932;
  wire  T_3933;
  wire  T_3934;
  wire  T_3935;
  wire  T_3936;
  wire  T_3937;
  wire [7:0] GEN_603;
  wire [8:0] T_3939;
  wire [7:0] T_3940;
  wire [7:0] GEN_604;
  wire [8:0] T_3942;
  wire [7:0] T_3943;
  wire [7:0] GEN_605;
  wire [8:0] T_3945;
  wire [7:0] T_3946;
  wire [7:0] GEN_606;
  wire [8:0] T_3948;
  wire [7:0] T_3949;
  wire [7:0] GEN_607;
  wire [8:0] T_3951;
  wire [7:0] T_3952;
  wire [7:0] GEN_608;
  wire [8:0] T_3954;
  wire [7:0] T_3955;
  wire [7:0] GEN_609;
  wire [8:0] T_3957;
  wire [7:0] T_3958;
  wire [7:0] GEN_610;
  wire [8:0] T_3960;
  wire [7:0] T_3961;
  wire [7:0] T_3967_0;
  wire [7:0] T_3967_1;
  wire [7:0] T_3967_2;
  wire [7:0] T_3967_3;
  wire [7:0] T_3967_4;
  wire [7:0] T_3967_5;
  wire [7:0] T_3967_6;
  wire [7:0] T_3967_7;
  wire [15:0] T_3969;
  wire [15:0] T_3970;
  wire [31:0] T_3971;
  wire [15:0] T_3972;
  wire [15:0] T_3973;
  wire [31:0] T_3974;
  wire [63:0] T_3975;
  wire [63:0] T_3976;
  wire [63:0] GEN_24;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [63:0] GEN_366;
  wire [63:0] GEN_367;
  wire [63:0] GEN_368;
  wire [63:0] GEN_369;
  wire [63:0] T_3977;
  wire [63:0] T_3978;
  wire [63:0] T_3979;
  wire [63:0] GEN_25;
  wire [63:0] GEN_370;
  wire [63:0] GEN_371;
  wire [63:0] GEN_372;
  wire [63:0] GEN_373;
  wire [63:0] GEN_374;
  wire [63:0] GEN_375;
  wire [63:0] GEN_376;
  wire [63:0] GEN_377;
  wire [7:0] T_3993_0;
  wire [7:0] T_4005;
  wire [7:0] GEN_26;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [7:0] GEN_381;
  wire [7:0] GEN_382;
  wire [7:0] GEN_383;
  wire [7:0] GEN_384;
  wire [7:0] T_4006;
  wire [7:0] GEN_27;
  wire [7:0] GEN_385;
  wire [7:0] GEN_386;
  wire [7:0] GEN_387;
  wire [7:0] GEN_388;
  wire [7:0] GEN_389;
  wire [7:0] GEN_390;
  wire [7:0] GEN_391;
  wire [7:0] GEN_392;
  wire [63:0] GEN_404;
  wire [63:0] GEN_405;
  wire [63:0] GEN_406;
  wire [63:0] GEN_407;
  wire [63:0] GEN_408;
  wire [63:0] GEN_409;
  wire [63:0] GEN_410;
  wire [63:0] GEN_411;
  wire [7:0] GEN_415;
  wire [7:0] GEN_416;
  wire [7:0] GEN_417;
  wire [7:0] GEN_418;
  wire [7:0] GEN_419;
  wire [7:0] GEN_420;
  wire [7:0] GEN_421;
  wire [7:0] GEN_422;
  wire  T_4009;
  wire  T_4010;
  wire  T_4011;
  wire  T_4012;
  wire  T_4013;
  wire  T_4014;
  wire  T_4015;
  wire  T_4017;
  wire  T_4019;
  wire [3:0] GEN_423;
  wire [7:0] GEN_424;
  wire [7:0] GEN_425;
  wire [7:0] GEN_426;
  wire [7:0] GEN_427;
  wire [7:0] GEN_428;
  wire [7:0] GEN_429;
  wire [7:0] GEN_430;
  wire [7:0] GEN_431;
  reg  GEN_28;
  reg [31:0] GEN_114;
  reg  GEN_29;
  reg [31:0] GEN_115;
  Queue_11 Queue_12_1 (
    .clk(Queue_12_1_clk),
    .reset(Queue_12_1_reset),
    .io_enq_ready(Queue_12_1_io_enq_ready),
    .io_enq_valid(Queue_12_1_io_enq_valid),
    .io_enq_bits_client_xact_id(Queue_12_1_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(Queue_12_1_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(Queue_12_1_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(Queue_12_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(Queue_12_1_io_enq_bits_a_type),
    .io_deq_ready(Queue_12_1_io_deq_ready),
    .io_deq_valid(Queue_12_1_io_deq_valid),
    .io_deq_bits_client_xact_id(Queue_12_1_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(Queue_12_1_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(Queue_12_1_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(Queue_12_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(Queue_12_1_io_deq_bits_a_type),
    .io_count(Queue_12_1_io_count)
  );
  assign io_inner_acquire_ready = T_2099;
  assign io_inner_grant_valid = GEN_361;
  assign io_inner_grant_bits_addr_beat = GEN_350;
  assign io_inner_grant_bits_client_xact_id = GEN_351;
  assign io_inner_grant_bits_manager_xact_id = GEN_352;
  assign io_inner_grant_bits_is_builtin_type = GEN_353;
  assign io_inner_grant_bits_g_type = GEN_354;
  assign io_inner_grant_bits_data = GEN_355;
  assign io_inner_grant_bits_client_id = GEN_356;
  assign io_inner_finish_ready = T_2977;
  assign io_inner_probe_valid = T_2211;
  assign io_inner_probe_bits_addr_block = T_2155_addr_block;
  assign io_inner_probe_bits_p_type = T_2155_p_type;
  assign io_inner_probe_bits_client_id = T_2155_client_id;
  assign io_inner_release_ready = T_2709;
  assign io_outer_acquire_valid = T_3169;
  assign io_outer_acquire_bits_addr_block = T_3369_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3369_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3369_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3369_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3369_a_type;
  assign io_outer_acquire_bits_union = T_3369_union;
  assign io_outer_acquire_bits_data = T_3369_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2996;
  assign io_outer_release_bits_addr_beat = T_3045_addr_beat;
  assign io_outer_release_bits_addr_block = T_3045_addr_block;
  assign io_outer_release_bits_client_xact_id = T_3045_client_xact_id;
  assign io_outer_release_bits_voluntary = T_3045_voluntary;
  assign io_outer_release_bits_r_type = T_3045_r_type;
  assign io_outer_release_bits_data = T_3045_data;
  assign io_outer_grant_ready = T_2977;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_28;
  assign io_outer_finish_bits_manager_id = GEN_29;
  assign io_alloc_iacq_matches = T_1842;
  assign io_alloc_iacq_can = T_1733;
  assign io_alloc_irel_matches = T_1845;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1848;
  assign io_alloc_oprb_can = 1'h0;
  assign T_44 = T_4017;
  assign T_69 = T_99_addr_beat;
  assign T_99_client_xact_id = T_1930_client_xact_id;
  assign T_99_addr_beat = T_1930_addr_beat;
  assign T_99_client_id = T_1930_client_id;
  assign T_99_is_builtin_type = T_1930_is_builtin_type;
  assign T_99_a_type = T_1930_a_type;
  assign T_144_pending = T_2380;
  assign T_144_up_idx = T_2319;
  assign T_144_up_done = T_2320;
  assign T_144_down_idx = T_2363;
  assign T_144_down_done = T_2364;
  assign T_153 = T_1960;
  assign T_155 = T_3808;
  assign T_157 = T_3809;
  assign T_166_pending = T_3559;
  assign T_166_up_idx = T_3527;
  assign T_166_up_done = T_3528;
  assign T_166_down_idx = 3'h0;
  assign T_166_down_done = T_3529;
  assign T_186_pending = T_3161;
  assign T_186_up_idx = T_3102;
  assign T_186_up_done = T_3103;
  assign T_186_down_idx = T_3144;
  assign T_186_down_done = T_3145;
  assign T_210_pending = T_2976;
  assign T_210_up_idx = T_2919;
  assign T_210_up_done = T_2920;
  assign T_210_down_idx = T_2959;
  assign T_210_down_done = T_2960;
  assign GEN_432 = {{7'd0}, 1'h0};
  assign T_219 = T_201 != GEN_432;
  assign T_220 = T_199 | T_219;
  assign T_221 = T_220 | T_210_pending;
  assign T_247_sharers = 1'h0;
  assign T_299_state = {{1'd0}, 1'h0};
  assign T_395_inner_sharers = T_247_sharers;
  assign T_395_outer_state = T_299_state;
  assign T_1733 = T_55 == 4'h0;
  assign T_1734 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1735 = T_1733 & T_1734;
  assign T_1736 = T_1735 & io_alloc_iacq_should;
  assign T_1745_0 = 3'h3;
  assign T_1747 = T_1745_0 == io_inner_acquire_bits_a_type;
  assign T_1750 = io_inner_acquire_bits_is_builtin_type & T_1747;
  assign T_1751 = T_1736 & T_1750;
  assign T_1760_0 = 3'h3;
  assign T_1762 = T_1760_0 == io_inner_acquire_bits_a_type;
  assign T_1765 = io_inner_acquire_bits_is_builtin_type & T_1762;
  assign T_1767 = T_1765 == 1'h0;
  assign GEN_433 = {{2'd0}, 1'h0};
  assign T_1769 = io_inner_acquire_bits_addr_beat == GEN_433;
  assign T_1770 = T_1767 | T_1769;
  assign T_1772 = T_1770 == 1'h0;
  assign T_1773 = T_1751 & T_1772;
  assign T_1775 = T_1773 == 1'h0;
  assign T_1776 = T_1775 | reset;
  assign T_1778 = T_1776 == 1'h0;
  assign T_1779 = T_55 != 4'h0;
  assign T_1780 = T_1779 & T_153;
  assign T_1782 = T_99_a_type == 3'h5;
  assign T_1784 = T_99_a_type == 3'h6;
  assign T_1785 = T_1782 | T_1784;
  assign T_1786 = T_99_is_builtin_type & T_1785;
  assign T_1787 = T_1780 & T_1786;
  assign T_1789 = T_1787 == 1'h0;
  assign T_1790 = T_1789 | reset;
  assign T_1792 = T_1790 == 1'h0;
  assign T_1796 = T_99_a_type == 3'h4;
  assign T_1797 = T_99_is_builtin_type & T_1796;
  assign T_1798 = T_1780 & T_1797;
  assign T_1800 = T_1798 == 1'h0;
  assign T_1801 = T_1800 | reset;
  assign T_1803 = T_1801 == 1'h0;
  assign T_1817_0 = 64'h0;
  assign T_1817_1 = 64'h0;
  assign T_1817_2 = 64'h0;
  assign T_1817_3 = 64'h0;
  assign T_1817_4 = 64'h0;
  assign T_1817_5 = 64'h0;
  assign T_1817_6 = 64'h0;
  assign T_1817_7 = 64'h0;
  assign T_1835_0 = 8'h0;
  assign T_1835_1 = 8'h0;
  assign T_1835_2 = 8'h0;
  assign T_1835_3 = 8'h0;
  assign T_1835_4 = 8'h0;
  assign T_1835_5 = 8'h0;
  assign T_1835_6 = 8'h0;
  assign T_1835_7 = 8'h0;
  assign T_1841 = io_inner_acquire_bits_addr_block == T_57;
  assign T_1842 = T_1779 & T_1841;
  assign T_1844 = io_inner_release_bits_addr_block == T_57;
  assign T_1845 = T_1779 & T_1844;
  assign T_1847 = io_outer_probe_bits_addr_block == T_57;
  assign T_1848 = T_1779 & T_1847;
  assign Queue_12_1_clk = clk;
  assign Queue_12_1_reset = reset;
  assign Queue_12_1_io_enq_valid = T_1929;
  assign Queue_12_1_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign Queue_12_1_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign Queue_12_1_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign Queue_12_1_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign Queue_12_1_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign Queue_12_1_io_deq_ready = GEN_349;
  assign T_1884 = T_1733 & io_alloc_iacq_should;
  assign T_1885 = T_1884 & io_inner_acquire_valid;
  assign T_1887 = T_99_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1896_0 = 3'h3;
  assign T_1898 = T_1896_0 == T_99_a_type;
  assign T_1901 = T_99_is_builtin_type & T_1898;
  assign T_1902 = T_1887 & T_1901;
  assign T_1903 = T_1902 & T_153;
  assign T_1904 = T_175 >> io_inner_acquire_bits_addr_beat;
  assign T_1905 = T_1904[0];
  assign T_1906 = T_1903 & T_1905;
  assign T_1908 = T_1906 & io_inner_acquire_valid;
  assign T_1917_0 = 3'h3;
  assign T_1919 = T_1917_0 == io_inner_acquire_bits_a_type;
  assign T_1922 = io_inner_acquire_bits_is_builtin_type & T_1919;
  assign T_1924 = T_1922 == 1'h0;
  assign T_1927 = T_1924 | T_1769;
  assign T_1928 = T_1908 & T_1927;
  assign T_1929 = T_1885 | T_1928;
  assign T_1930_client_xact_id = Queue_12_1_io_deq_valid ? Queue_12_1_io_deq_bits_client_xact_id : Queue_12_1_io_enq_bits_client_xact_id;
  assign T_1930_addr_beat = Queue_12_1_io_deq_valid ? Queue_12_1_io_deq_bits_addr_beat : Queue_12_1_io_enq_bits_addr_beat;
  assign T_1930_client_id = Queue_12_1_io_deq_valid ? Queue_12_1_io_deq_bits_client_id : Queue_12_1_io_enq_bits_client_id;
  assign T_1930_is_builtin_type = Queue_12_1_io_deq_valid ? Queue_12_1_io_deq_bits_is_builtin_type : Queue_12_1_io_enq_bits_is_builtin_type;
  assign T_1930_a_type = Queue_12_1_io_deq_valid ? Queue_12_1_io_deq_bits_a_type : Queue_12_1_io_enq_bits_a_type;
  assign GEN_435 = {{1'd0}, 1'h0};
  assign T_1960 = Queue_12_1_io_count > GEN_435;
  assign T_1962 = T_1779 | io_alloc_iacq_should;
  assign T_1972_0 = 3'h2;
  assign T_1972_1 = 3'h3;
  assign T_1972_2 = 3'h4;
  assign T_1974 = T_1972_0 == io_inner_acquire_bits_a_type;
  assign T_1975 = T_1972_1 == io_inner_acquire_bits_a_type;
  assign T_1976 = T_1972_2 == io_inner_acquire_bits_a_type;
  assign T_1979 = T_1974 | T_1975;
  assign T_1980 = T_1979 | T_1976;
  assign T_1981 = io_inner_acquire_bits_is_builtin_type & T_1980;
  assign T_1982 = T_1734 & T_1981;
  assign GEN_436 = {{7'd0}, T_1982};
  assign T_1984 = 8'h0 - GEN_436;
  assign T_1985 = T_1984[7:0];
  assign T_1986 = ~ T_1985;
  assign GEN_437 = {{7'd0}, 1'h1};
  assign T_1988 = GEN_437 << io_inner_acquire_bits_addr_beat;
  assign T_1989 = ~ T_1988;
  assign T_1990 = T_1986 | T_1989;
  assign T_1991 = T_175 & T_1990;
  assign T_2001_0 = 3'h3;
  assign T_2003 = T_2001_0 == io_inner_acquire_bits_a_type;
  assign T_2006 = io_inner_acquire_bits_is_builtin_type & T_2003;
  assign T_2007 = T_1734 & T_2006;
  assign T_2010 = T_2007 & T_1769;
  assign T_2019 = T_2010 ? 8'hfe : 8'h0;
  assign T_2020 = T_1991 | T_2019;
  assign GEN_32 = T_1962 ? T_2020 : T_175;
  assign GEN_439 = {{3'd0}, 1'h0};
  assign T_2028 = 4'h8 * GEN_439;
  assign T_2030 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_2031 = io_inner_acquire_bits_is_builtin_type & T_2030;
  assign T_2033 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_2034 = io_inner_acquire_bits_is_builtin_type & T_2033;
  assign T_2035 = T_2031 | T_2034;
  assign T_2036 = io_inner_acquire_bits_union[5:1];
  assign T_2037 = T_2035 ? 5'h1 : T_2036;
  assign T_2038 = io_inner_acquire_bits_union[11:9];
  assign T_2039 = io_inner_acquire_bits_union[8:6];
  assign T_2052_0 = 3'h2;
  assign T_2052_1 = 3'h3;
  assign T_2052_2 = 3'h4;
  assign T_2054 = T_2052_0 == io_inner_acquire_bits_a_type;
  assign T_2055 = T_2052_1 == io_inner_acquire_bits_a_type;
  assign T_2056 = T_2052_2 == io_inner_acquire_bits_a_type;
  assign T_2059 = T_2054 | T_2055;
  assign T_2060 = T_2059 | T_2056;
  assign T_2061 = io_inner_acquire_bits_is_builtin_type & T_2060;
  assign T_2062 = T_1734 & T_2061;
  assign GEN_440 = {{7'd0}, T_2062};
  assign T_2064 = 8'h0 - GEN_440;
  assign T_2065 = T_2064[7:0];
  assign T_2066 = ~ T_2065;
  assign T_2070 = T_2066 | T_1989;
  assign T_2072 = T_2034 ? T_2070 : {{7'd0}, 1'h0};
  assign GEN_33 = T_1885 ? io_inner_acquire_bits_addr_block : T_57;
  assign GEN_34 = T_1885 ? 1'h0 : T_59;
  assign GEN_35 = T_1885 ? T_2028 : T_61;
  assign GEN_36 = T_1885 ? T_2037 : T_63;
  assign GEN_37 = T_1885 ? T_2038 : T_65;
  assign GEN_38 = T_1885 ? T_2039 : T_67;
  assign GEN_42 = T_1885 ? T_2072 : GEN_32;
  assign GEN_43 = T_1885 ? {{7'd0}, 1'h0} : T_177;
  assign GEN_44 = T_1885 ? 4'h5 : T_55;
  assign T_2075 = T_175 != GEN_432;
  assign T_2088_0 = 3'h3;
  assign T_2090 = T_2088_0 == T_99_a_type;
  assign T_2093 = T_99_is_builtin_type & T_2090;
  assign T_2094 = T_1887 & T_2093;
  assign T_2095 = T_2094 & T_153;
  assign T_2098 = T_2095 & T_1905;
  assign T_2099 = T_1733 | T_2098;
  assign T_2100 = ~ T_177;
  assign skip_outer_acquire = T_2100 == GEN_432;
  assign T_2109 = 3'h4 == T_99_a_type;
  assign T_2110 = T_2109 ? 2'h0 : 2'h2;
  assign T_2111 = 3'h6 == T_99_a_type;
  assign T_2112 = T_2111 ? 2'h0 : T_2110;
  assign T_2113 = 3'h5 == T_99_a_type;
  assign T_2114 = T_2113 ? 2'h2 : T_2112;
  assign T_2115 = 3'h2 == T_99_a_type;
  assign T_2116 = T_2115 ? 2'h0 : T_2114;
  assign T_2117 = 3'h0 == T_99_a_type;
  assign T_2118 = T_2117 ? 2'h2 : T_2116;
  assign T_2119 = 3'h3 == T_99_a_type;
  assign T_2120 = T_2119 ? 2'h0 : T_2118;
  assign T_2121 = 3'h1 == T_99_a_type;
  assign T_2122 = T_2121 ? 2'h2 : T_2120;
  assign GEN_444 = {{2'd0}, 1'h1};
  assign T_2123 = GEN_444 == T_99_a_type;
  assign T_2124 = T_2123 ? 2'h0 : 2'h2;
  assign T_2125 = GEN_433 == T_99_a_type;
  assign T_2126 = T_2125 ? 2'h1 : T_2124;
  assign T_2127 = T_99_is_builtin_type ? T_2122 : T_2126;
  assign T_2155_addr_block = T_57;
  assign T_2155_p_type = T_2127;
  assign T_2155_client_id = 1'h0;
  assign T_2183 = skip_outer_acquire == 1'h0;
  assign T_2184 = T_2183 ? 4'h6 : 4'h7;
  assign T_2193_pending = T_2276;
  assign T_2193_up_idx = 3'h0;
  assign T_2193_up_done = T_2201;
  assign T_2193_down_idx = T_2259;
  assign T_2193_down_done = T_2260;
  assign T_2201 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2202 = ~ T_2201;
  assign GEN_446 = {{1'd0}, 1'h1};
  assign T_2204 = GEN_446 << io_inner_probe_bits_client_id;
  assign T_2205 = ~ T_2204;
  assign GEN_447 = {{1'd0}, T_2202};
  assign T_2206 = GEN_447 | T_2205;
  assign GEN_448 = {{1'd0}, T_195};
  assign T_2207 = GEN_448 & T_2206;
  assign T_2208 = T_55 == 4'h5;
  assign T_2211 = T_2208 & T_195;
  assign T_2228 = io_inner_release_ready & io_inner_release_valid;
  assign T_2231 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2232 = T_1779 & T_2231;
  assign T_2233 = T_2228 & T_2232;
  assign T_2240_0 = 3'h0;
  assign T_2240_1 = 3'h1;
  assign T_2240_2 = 3'h2;
  assign T_2242 = T_2240_0 == io_inner_release_bits_r_type;
  assign T_2243 = T_2240_1 == io_inner_release_bits_r_type;
  assign T_2244 = T_2240_2 == io_inner_release_bits_r_type;
  assign T_2247 = T_2242 | T_2243;
  assign T_2248 = T_2247 | T_2244;
  assign T_2250 = T_2233 & T_2248;
  assign T_2254 = T_2252 == 3'h7;
  assign T_2256 = T_2252 + GEN_444;
  assign T_2257 = T_2256[2:0];
  assign GEN_46 = T_2250 ? T_2257 : T_2252;
  assign T_2258 = T_2250 & T_2254;
  assign T_2259 = T_2248 ? T_2252 : {{2'd0}, 1'h0};
  assign T_2260 = T_2248 ? T_2258 : T_2233;
  assign T_2264 = T_2260 == 1'h0;
  assign T_2265 = T_2201 & T_2264;
  assign T_2267 = T_2262 + 1'h1;
  assign T_2268 = T_2267[0:0];
  assign GEN_47 = T_2265 ? T_2268 : T_2262;
  assign T_2270 = T_2201 == 1'h0;
  assign T_2271 = T_2260 & T_2270;
  assign T_2273 = T_2262 - 1'h1;
  assign T_2274 = T_2273[0:0];
  assign GEN_48 = T_2271 ? T_2274 : GEN_47;
  assign T_2276 = T_2262 > 1'h0;
  assign T_2280 = T_195 | T_2193_pending;
  assign T_2282 = T_2280 == 1'h0;
  assign T_2283 = T_2208 & T_2282;
  assign GEN_49 = T_2283 ? T_2184 : GEN_44;
  assign T_2287 = T_1733 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2288 = T_2287 & io_inner_release_bits_voluntary;
  assign T_2293 = T_2228 & T_2288;
  assign T_2300_0 = 3'h0;
  assign T_2300_1 = 3'h1;
  assign T_2300_2 = 3'h2;
  assign T_2302 = T_2300_0 == io_inner_release_bits_r_type;
  assign T_2303 = T_2300_1 == io_inner_release_bits_r_type;
  assign T_2304 = T_2300_2 == io_inner_release_bits_r_type;
  assign T_2307 = T_2302 | T_2303;
  assign T_2308 = T_2307 | T_2304;
  assign T_2310 = T_2293 & T_2308;
  assign T_2314 = T_2312 == 3'h7;
  assign T_2316 = T_2312 + GEN_444;
  assign T_2317 = T_2316[2:0];
  assign GEN_50 = T_2310 ? T_2317 : T_2312;
  assign T_2318 = T_2310 & T_2314;
  assign T_2319 = T_2308 ? T_2312 : {{2'd0}, 1'h0};
  assign T_2320 = T_2308 ? T_2318 : T_2293;
  assign T_2321 = io_inner_grant_ready & io_inner_grant_valid;
  assign GEN_452 = {{1'd0}, 3'h0};
  assign T_2324 = io_inner_grant_bits_g_type == GEN_452;
  assign T_2325 = io_inner_grant_bits_is_builtin_type & T_2324;
  assign T_2326 = T_1779 & T_2325;
  assign T_2327 = T_2321 & T_2326;
  assign T_2335_0 = 3'h5;
  assign GEN_453 = {{1'd0}, T_2335_0};
  assign T_2337 = GEN_453 == io_inner_grant_bits_g_type;
  assign T_2345_0 = 2'h0;
  assign T_2345_1 = 2'h1;
  assign GEN_454 = {{2'd0}, T_2345_0};
  assign T_2347 = GEN_454 == io_inner_grant_bits_g_type;
  assign GEN_455 = {{2'd0}, T_2345_1};
  assign T_2348 = GEN_455 == io_inner_grant_bits_g_type;
  assign T_2351 = T_2347 | T_2348;
  assign T_2352 = io_inner_grant_bits_is_builtin_type ? T_2337 : T_2351;
  assign T_2354 = T_2327 & T_2352;
  assign T_2358 = T_2356 == 3'h7;
  assign T_2360 = T_2356 + GEN_444;
  assign T_2361 = T_2360[2:0];
  assign GEN_51 = T_2354 ? T_2361 : T_2356;
  assign T_2362 = T_2354 & T_2358;
  assign T_2363 = T_2352 ? T_2356 : {{2'd0}, 1'h0};
  assign T_2364 = T_2352 ? T_2362 : T_2327;
  assign T_2368 = T_2364 == 1'h0;
  assign T_2369 = T_2320 & T_2368;
  assign T_2371 = T_2366 + 1'h1;
  assign T_2372 = T_2371[0:0];
  assign GEN_52 = T_2369 ? T_2372 : T_2366;
  assign T_2374 = T_2320 == 1'h0;
  assign T_2375 = T_2364 & T_2374;
  assign T_2377 = T_2366 - 1'h1;
  assign T_2378 = T_2377[0:0];
  assign GEN_53 = T_2375 ? T_2378 : GEN_52;
  assign T_2380 = T_2366 > 1'h0;
  assign T_2382 = T_1733 & io_alloc_irel_should;
  assign T_2383 = T_2382 & io_inner_release_valid;
  assign GEN_54 = T_2383 ? io_inner_release_bits_addr_block : GEN_33;
  assign GEN_55 = T_2383 ? 4'h7 : GEN_49;
  assign T_2386 = T_1844 & io_inner_release_bits_voluntary;
  assign T_2392_0 = 4'h0;
  assign T_2392_1 = 4'h8;
  assign T_2394 = T_2392_0 == T_55;
  assign T_2395 = T_2392_1 == T_55;
  assign T_2398 = T_2394 | T_2395;
  assign T_2400 = T_2398 == 1'h0;
  assign T_2401 = T_2386 & T_2400;
  assign T_2403 = T_44 == 1'h0;
  assign T_2404 = T_2401 & T_2403;
  assign T_2405 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2407 = T_2405 == 1'h0;
  assign T_2408 = T_2404 & T_2407;
  assign T_2411 = T_2321 == 1'h0;
  assign T_2412 = T_2408 & T_2411;
  assign T_2414 = T_144_pending == 1'h0;
  assign T_2415 = T_2412 & T_2414;
  assign T_2422_0 = 3'h0;
  assign T_2422_1 = 3'h1;
  assign T_2422_2 = 3'h2;
  assign T_2424 = T_2422_0 == io_inner_release_bits_r_type;
  assign T_2425 = T_2422_1 == io_inner_release_bits_r_type;
  assign T_2426 = T_2422_2 == io_inner_release_bits_r_type;
  assign T_2429 = T_2424 | T_2425;
  assign T_2430 = T_2429 | T_2426;
  assign T_2433 = T_2430 == 1'h0;
  assign T_2435 = io_inner_release_bits_addr_beat == GEN_433;
  assign T_2436 = T_2433 | T_2435;
  assign T_2437 = T_2415 & T_2436;
  assign T_2438 = io_alloc_irel_should | T_2437;
  assign T_2445_0 = 3'h0;
  assign T_2445_1 = 3'h1;
  assign T_2445_2 = 3'h2;
  assign T_2447 = T_2445_0 == io_inner_release_bits_r_type;
  assign T_2448 = T_2445_1 == io_inner_release_bits_r_type;
  assign T_2449 = T_2445_2 == io_inner_release_bits_r_type;
  assign T_2452 = T_2447 | T_2448;
  assign T_2453 = T_2452 | T_2449;
  assign T_2461_0 = 3'h0;
  assign T_2461_1 = 3'h1;
  assign T_2461_2 = 3'h2;
  assign T_2463 = T_2461_0 == io_inner_release_bits_r_type;
  assign T_2464 = T_2461_1 == io_inner_release_bits_r_type;
  assign T_2465 = T_2461_2 == io_inner_release_bits_r_type;
  assign T_2468 = T_2463 | T_2464;
  assign T_2469 = T_2468 | T_2465;
  assign T_2470 = T_2228 & T_2469;
  assign GEN_458 = {{7'd0}, T_2470};
  assign T_2472 = 8'h0 - GEN_458;
  assign T_2473 = T_2472[7:0];
  assign T_2474 = ~ T_2473;
  assign T_2476 = GEN_437 << io_inner_release_bits_addr_beat;
  assign T_2477 = ~ T_2476;
  assign T_2478 = T_2474 | T_2477;
  assign T_2480 = T_2453 ? T_2478 : {{7'd0}, 1'h0};
  assign GEN_56 = T_2438 ? io_inner_release_bits_r_type : T_129;
  assign GEN_57 = T_2438 ? io_inner_release_bits_client_id : T_131;
  assign GEN_58 = T_2438 ? io_inner_release_bits_client_xact_id : T_133;
  assign GEN_65 = T_2438 ? T_2480 : T_135;
  assign T_2484 = T_1844 & T_2231;
  assign T_2486 = T_2484 & T_2208;
  assign T_2488 = T_2438 == 1'h0;
  assign T_2489 = T_2488 & T_2486;
  assign T_2496_0 = 3'h0;
  assign T_2496_1 = 3'h1;
  assign T_2496_2 = 3'h2;
  assign T_2498 = T_2496_0 == io_inner_release_bits_r_type;
  assign T_2499 = T_2496_1 == io_inner_release_bits_r_type;
  assign T_2500 = T_2496_2 == io_inner_release_bits_r_type;
  assign T_2503 = T_2498 | T_2499;
  assign T_2504 = T_2503 | T_2500;
  assign T_2505 = T_2228 & T_2504;
  assign GEN_460 = {{7'd0}, T_2505};
  assign T_2507 = 8'h0 - GEN_460;
  assign T_2508 = T_2507[7:0];
  assign T_2509 = ~ T_2508;
  assign T_2513 = T_2509 | T_2477;
  assign T_2514 = T_135 & T_2513;
  assign GEN_69 = T_2489 ? T_2514 : GEN_65;
  assign GEN_75 = T_2228 ? GEN_56 : T_129;
  assign GEN_76 = T_2228 ? GEN_57 : T_131;
  assign GEN_77 = T_2228 ? GEN_58 : T_133;
  assign GEN_84 = T_2228 ? GEN_69 : T_135;
  assign T_2520_0 = 4'h3;
  assign T_2520_1 = 4'h4;
  assign T_2520_2 = 4'h5;
  assign T_2520_3 = 4'h7;
  assign T_2522 = T_2520_0 == T_55;
  assign T_2523 = T_2520_1 == T_55;
  assign T_2524 = T_2520_2 == T_55;
  assign T_2525 = T_2520_3 == T_55;
  assign T_2528 = T_2522 | T_2523;
  assign T_2529 = T_2528 | T_2524;
  assign T_2530 = T_2529 | T_2525;
  assign T_2531 = T_2530 & T_144_pending;
  assign T_2533 = T_135 != GEN_432;
  assign T_2534 = T_2533 | T_210_pending;
  assign T_2536 = T_2534 == 1'h0;
  assign T_2537 = T_2531 & T_2536;
  assign T_2572_addr_beat = {{2'd0}, 1'h0};
  assign T_2572_addr_block = T_57;
  assign T_2572_client_xact_id = T_133;
  assign T_2572_voluntary = 1'h1;
  assign T_2572_r_type = T_129;
  assign T_2572_data = {{63'd0}, 1'h0};
  assign T_2572_client_id = T_131;
  assign T_2639_addr_beat = {{2'd0}, 1'h0};
  assign T_2639_client_xact_id = T_2572_client_xact_id;
  assign T_2639_manager_xact_id = {{2'd0}, 1'h0};
  assign T_2639_is_builtin_type = 1'h1;
  assign T_2639_g_type = {{1'd0}, 3'h0};
  assign T_2639_data = {{63'd0}, 1'h0};
  assign T_2639_client_id = T_2572_client_id;
  assign T_2679_0 = 4'h0;
  assign T_2679_1 = 4'h8;
  assign T_2681 = T_2679_0 == T_55;
  assign T_2682 = T_2679_1 == T_55;
  assign T_2685 = T_2681 | T_2682;
  assign T_2687 = T_2685 == 1'h0;
  assign T_2688 = T_2386 & T_2687;
  assign T_2691 = T_2688 & T_2403;
  assign T_2695 = T_2691 & T_2407;
  assign T_2699 = T_2695 & T_2411;
  assign T_2702 = T_2699 & T_2414;
  assign T_2709 = T_2702 | T_2486;
  assign T_2716_0 = 3'h0;
  assign T_2716_1 = 3'h1;
  assign T_2716_2 = 3'h2;
  assign T_2718 = T_2716_0 == io_inner_release_bits_r_type;
  assign T_2719 = T_2716_1 == io_inner_release_bits_r_type;
  assign T_2720 = T_2716_2 == io_inner_release_bits_r_type;
  assign T_2723 = T_2718 | T_2719;
  assign T_2724 = T_2723 | T_2720;
  assign T_2725 = T_2228 & T_2724;
  assign GEN_0 = GEN_94;
  assign GEN_88 = GEN_444 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_465 = {{1'd0}, 2'h2};
  assign GEN_89 = GEN_465 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_88;
  assign GEN_466 = {{1'd0}, 2'h3};
  assign GEN_90 = GEN_466 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_89;
  assign GEN_91 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_90;
  assign GEN_92 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_91;
  assign GEN_93 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_92;
  assign GEN_94 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_93;
  assign T_2726 = GEN_0[0];
  assign GEN_1 = GEN_94;
  assign T_2727 = GEN_1[1];
  assign GEN_2 = GEN_94;
  assign T_2728 = GEN_2[2];
  assign GEN_3 = GEN_94;
  assign T_2729 = GEN_3[3];
  assign GEN_4 = GEN_94;
  assign T_2730 = GEN_4[4];
  assign GEN_5 = GEN_94;
  assign T_2731 = GEN_5[5];
  assign GEN_6 = GEN_94;
  assign T_2732 = GEN_6[6];
  assign GEN_7 = GEN_94;
  assign T_2733 = GEN_7[7];
  assign GEN_488 = {{7'd0}, T_2726};
  assign T_2735 = 8'h0 - GEN_488;
  assign T_2736 = T_2735[7:0];
  assign GEN_489 = {{7'd0}, T_2727};
  assign T_2738 = 8'h0 - GEN_489;
  assign T_2739 = T_2738[7:0];
  assign GEN_490 = {{7'd0}, T_2728};
  assign T_2741 = 8'h0 - GEN_490;
  assign T_2742 = T_2741[7:0];
  assign GEN_491 = {{7'd0}, T_2729};
  assign T_2744 = 8'h0 - GEN_491;
  assign T_2745 = T_2744[7:0];
  assign GEN_492 = {{7'd0}, T_2730};
  assign T_2747 = 8'h0 - GEN_492;
  assign T_2748 = T_2747[7:0];
  assign GEN_493 = {{7'd0}, T_2731};
  assign T_2750 = 8'h0 - GEN_493;
  assign T_2751 = T_2750[7:0];
  assign GEN_494 = {{7'd0}, T_2732};
  assign T_2753 = 8'h0 - GEN_494;
  assign T_2754 = T_2753[7:0];
  assign GEN_495 = {{7'd0}, T_2733};
  assign T_2756 = 8'h0 - GEN_495;
  assign T_2757 = T_2756[7:0];
  assign T_2763_0 = T_2736;
  assign T_2763_1 = T_2739;
  assign T_2763_2 = T_2742;
  assign T_2763_3 = T_2745;
  assign T_2763_4 = T_2748;
  assign T_2763_5 = T_2751;
  assign T_2763_6 = T_2754;
  assign T_2763_7 = T_2757;
  assign T_2765 = {T_2763_1,T_2763_0};
  assign T_2766 = {T_2763_3,T_2763_2};
  assign T_2767 = {T_2766,T_2765};
  assign T_2768 = {T_2763_5,T_2763_4};
  assign T_2769 = {T_2763_7,T_2763_6};
  assign T_2770 = {T_2769,T_2768};
  assign T_2771 = {T_2770,T_2767};
  assign T_2772 = ~ T_2771;
  assign T_2773 = T_2772 & io_inner_release_bits_data;
  assign GEN_8 = GEN_150;
  assign GEN_144 = GEN_444 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_145 = GEN_465 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_144;
  assign GEN_146 = GEN_466 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_145;
  assign GEN_147 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_146;
  assign GEN_148 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_147;
  assign GEN_149 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_148;
  assign GEN_150 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_149;
  assign T_2774 = T_2771 & GEN_8;
  assign T_2775 = T_2773 | T_2774;
  assign GEN_9 = T_2775;
  assign GEN_151 = GEN_433 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_152 = GEN_444 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_153 = GEN_465 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_154 = GEN_466 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_155 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_156 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_157 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_158 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_177 = T_2725 ? GEN_151 : data_buffer_0;
  assign GEN_178 = T_2725 ? GEN_152 : data_buffer_1;
  assign GEN_179 = T_2725 ? GEN_153 : data_buffer_2;
  assign GEN_180 = T_2725 ? GEN_154 : data_buffer_3;
  assign GEN_181 = T_2725 ? GEN_155 : data_buffer_4;
  assign GEN_182 = T_2725 ? GEN_156 : data_buffer_5;
  assign GEN_183 = T_2725 ? GEN_157 : data_buffer_6;
  assign GEN_184 = T_2725 ? GEN_158 : data_buffer_7;
  assign T_2806_state = 2'h2;
  assign T_2832 = T_1779 | io_alloc_irel_should;
  assign T_2833 = io_outer_release_ready & io_outer_release_valid;
  assign T_2839_0 = 3'h0;
  assign T_2839_1 = 3'h1;
  assign T_2839_2 = 3'h2;
  assign T_2841 = T_2839_0 == io_outer_release_bits_r_type;
  assign T_2842 = T_2839_1 == io_outer_release_bits_r_type;
  assign T_2843 = T_2839_2 == io_outer_release_bits_r_type;
  assign T_2846 = T_2841 | T_2842;
  assign T_2847 = T_2846 | T_2843;
  assign T_2848 = T_2833 & T_2847;
  assign GEN_503 = {{7'd0}, T_2848};
  assign T_2850 = 8'h0 - GEN_503;
  assign T_2851 = T_2850[7:0];
  assign T_2852 = ~ T_2851;
  assign T_2854 = GEN_437 << io_outer_release_bits_addr_beat;
  assign T_2855 = ~ T_2854;
  assign T_2856 = T_2852 | T_2855;
  assign T_2857 = T_201 & T_2856;
  assign T_2865_0 = 3'h0;
  assign T_2865_1 = 3'h1;
  assign T_2865_2 = 3'h2;
  assign T_2867 = T_2865_0 == io_inner_release_bits_r_type;
  assign T_2868 = T_2865_1 == io_inner_release_bits_r_type;
  assign T_2869 = T_2865_2 == io_inner_release_bits_r_type;
  assign T_2872 = T_2867 | T_2868;
  assign T_2873 = T_2872 | T_2869;
  assign T_2874 = T_2228 & T_2873;
  assign GEN_505 = {{7'd0}, T_2874};
  assign T_2877 = 8'h0 - GEN_505;
  assign T_2878 = T_2877[7:0];
  assign T_2881 = T_2878 & T_2476;
  assign T_2882 = T_2857 | T_2881;
  assign T_2883 = T_2882 | GEN_432;
  assign GEN_191 = T_2832 ? T_2883 : T_201;
  assign GEN_193 = T_2833 ? 1'h0 : T_199;
  assign T_2893 = T_2833 & io_outer_release_bits_voluntary;
  assign T_2900_0 = 3'h0;
  assign T_2900_1 = 3'h1;
  assign T_2900_2 = 3'h2;
  assign T_2902 = T_2900_0 == io_outer_release_bits_r_type;
  assign T_2903 = T_2900_1 == io_outer_release_bits_r_type;
  assign T_2904 = T_2900_2 == io_outer_release_bits_r_type;
  assign T_2907 = T_2902 | T_2903;
  assign T_2908 = T_2907 | T_2904;
  assign T_2910 = T_2893 & T_2908;
  assign T_2914 = T_2912 == 3'h7;
  assign T_2916 = T_2912 + GEN_444;
  assign T_2917 = T_2916[2:0];
  assign GEN_194 = T_2910 ? T_2917 : T_2912;
  assign T_2918 = T_2910 & T_2914;
  assign T_2919 = T_2908 ? T_2912 : {{2'd0}, 1'h0};
  assign T_2920 = T_2908 ? T_2918 : T_2893;
  assign T_2923 = io_outer_grant_bits_g_type == GEN_452;
  assign T_2924 = io_outer_grant_bits_is_builtin_type & T_2923;
  assign T_2925 = T_2405 & T_2924;
  assign T_2933_0 = 3'h5;
  assign GEN_510 = {{1'd0}, T_2933_0};
  assign T_2935 = GEN_510 == io_outer_grant_bits_g_type;
  assign T_2943_0 = 1'h0;
  assign GEN_511 = {{3'd0}, T_2943_0};
  assign T_2945 = GEN_511 == io_outer_grant_bits_g_type;
  assign T_2948 = io_outer_grant_bits_is_builtin_type ? T_2935 : T_2945;
  assign T_2950 = T_2925 & T_2948;
  assign T_2954 = T_2952 == 3'h7;
  assign T_2956 = T_2952 + GEN_444;
  assign T_2957 = T_2956[2:0];
  assign GEN_195 = T_2950 ? T_2957 : T_2952;
  assign T_2958 = T_2950 & T_2954;
  assign T_2959 = T_2948 ? T_2952 : {{2'd0}, 1'h0};
  assign T_2960 = T_2948 ? T_2958 : T_2925;
  assign T_2964 = T_2960 == 1'h0;
  assign T_2965 = T_2920 & T_2964;
  assign T_2967 = T_2962 + 1'h1;
  assign T_2968 = T_2967[0:0];
  assign GEN_196 = T_2965 ? T_2968 : T_2962;
  assign T_2970 = T_2920 == 1'h0;
  assign T_2971 = T_2960 & T_2970;
  assign T_2973 = T_2962 - 1'h1;
  assign T_2974 = T_2973[0:0];
  assign GEN_197 = T_2971 ? T_2974 : GEN_196;
  assign T_2976 = T_2962 > 1'h0;
  assign T_2977 = T_55 == 4'h7;
  assign T_2983_0 = 3'h0;
  assign T_2983_1 = 3'h1;
  assign T_2983_2 = 3'h2;
  assign T_2985 = T_2983_0 == io_outer_release_bits_r_type;
  assign T_2986 = T_2983_1 == io_outer_release_bits_r_type;
  assign T_2987 = T_2983_2 == io_outer_release_bits_r_type;
  assign T_2990 = T_2985 | T_2986;
  assign T_2991 = T_2990 | T_2987;
  assign T_2992 = T_201 >> T_210_up_idx;
  assign T_2993 = T_2992[0];
  assign T_2995 = T_2991 ? T_2993 : T_221;
  assign T_2996 = T_2977 & T_2995;
  assign T_3004_0 = 2'h2;
  assign T_3006 = T_3004_0 == T_2806_state;
  assign T_3009 = T_3006 ? 3'h0 : 3'h3;
  assign T_3045_addr_beat = T_210_up_idx;
  assign T_3045_addr_block = T_57;
  assign T_3045_client_xact_id = {{2'd0}, 1'h0};
  assign T_3045_voluntary = 1'h1;
  assign T_3045_r_type = T_3009;
  assign T_3045_data = GEN_10;
  assign GEN_10 = GEN_204;
  assign GEN_198 = GEN_444 == T_210_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_199 = GEN_465 == T_210_up_idx ? data_buffer_2 : GEN_198;
  assign GEN_200 = GEN_466 == T_210_up_idx ? data_buffer_3 : GEN_199;
  assign GEN_201 = 3'h4 == T_210_up_idx ? data_buffer_4 : GEN_200;
  assign GEN_202 = 3'h5 == T_210_up_idx ? data_buffer_5 : GEN_201;
  assign GEN_203 = 3'h6 == T_210_up_idx ? data_buffer_6 : GEN_202;
  assign GEN_204 = 3'h7 == T_210_up_idx ? data_buffer_7 : GEN_203;
  assign T_3074 = T_99_is_builtin_type == 1'h0;
  assign T_3076 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_3087_0 = 3'h3;
  assign T_3089 = T_3087_0 == io_outer_acquire_bits_a_type;
  assign T_3092 = io_outer_acquire_bits_is_builtin_type & T_3089;
  assign T_3093 = T_3076 & T_3092;
  assign T_3097 = T_3095 == 3'h7;
  assign T_3099 = T_3095 + GEN_444;
  assign T_3100 = T_3099[2:0];
  assign GEN_205 = T_3093 ? T_3100 : T_3095;
  assign T_3101 = T_3093 & T_3097;
  assign T_3102 = T_3092 ? T_3095 : T_69;
  assign T_3103 = T_3092 ? T_3101 : T_3076;
  assign T_3109 = T_2924 == 1'h0;
  assign T_3110 = T_2405 & T_3109;
  assign T_3118_0 = 3'h5;
  assign GEN_518 = {{1'd0}, T_3118_0};
  assign T_3120 = GEN_518 == io_outer_grant_bits_g_type;
  assign T_3128_0 = 1'h0;
  assign GEN_519 = {{3'd0}, T_3128_0};
  assign T_3130 = GEN_519 == io_outer_grant_bits_g_type;
  assign T_3133 = io_outer_grant_bits_is_builtin_type ? T_3120 : T_3130;
  assign T_3135 = T_3110 & T_3133;
  assign T_3139 = T_3137 == 3'h7;
  assign T_3141 = T_3137 + GEN_444;
  assign T_3142 = T_3141[2:0];
  assign GEN_206 = T_3135 ? T_3142 : T_3137;
  assign T_3143 = T_3135 & T_3139;
  assign T_3144 = T_3133 ? T_3137 : T_69;
  assign T_3145 = T_3133 ? T_3143 : T_3110;
  assign T_3149 = T_3145 == 1'h0;
  assign T_3150 = T_3103 & T_3149;
  assign T_3152 = T_3147 + 1'h1;
  assign T_3153 = T_3152[0:0];
  assign GEN_207 = T_3150 ? T_3153 : T_3147;
  assign T_3155 = T_3103 == 1'h0;
  assign T_3156 = T_3145 & T_3155;
  assign T_3158 = T_3147 - 1'h1;
  assign T_3159 = T_3158[0:0];
  assign GEN_208 = T_3156 ? T_3159 : GEN_207;
  assign T_3161 = T_3147 > 1'h0;
  assign T_3162 = T_55 == 4'h6;
  assign T_3163 = T_175 >> T_186_up_idx;
  assign T_3164 = T_3163[0];
  assign T_3166 = T_3164 == 1'h0;
  assign T_3168 = T_59 | T_3166;
  assign T_3169 = T_3162 & T_3168;
  assign T_3172 = T_63 == 5'h1;
  assign T_3173 = T_63 == 5'h7;
  assign T_3174 = T_3172 | T_3173;
  assign T_3175 = T_63[3];
  assign T_3176 = T_63 == 5'h4;
  assign T_3177 = T_3175 | T_3176;
  assign T_3178 = T_3174 | T_3177;
  assign T_3179 = T_63 == 5'h3;
  assign T_3180 = T_3178 | T_3179;
  assign T_3181 = T_63 == 5'h6;
  assign T_3182 = T_3180 | T_3181;
  assign T_3185 = {T_63,1'h1};
  assign T_3216_addr_block = T_57;
  assign T_3216_client_xact_id = {{2'd0}, 1'h0};
  assign T_3216_addr_beat = {{2'd0}, 1'h0};
  assign T_3216_is_builtin_type = 1'h0;
  assign T_3216_a_type = {{2'd0}, T_3182};
  assign T_3216_union = {{6'd0}, T_3185};
  assign T_3216_data = {{63'd0}, 1'h0};
  assign GEN_11 = GEN_215;
  assign GEN_209 = GEN_444 == T_186_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_210 = GEN_465 == T_186_up_idx ? wmask_buffer_2 : GEN_209;
  assign GEN_211 = GEN_466 == T_186_up_idx ? wmask_buffer_3 : GEN_210;
  assign GEN_212 = 3'h4 == T_186_up_idx ? wmask_buffer_4 : GEN_211;
  assign GEN_213 = 3'h5 == T_186_up_idx ? wmask_buffer_5 : GEN_212;
  assign GEN_214 = 3'h6 == T_186_up_idx ? wmask_buffer_6 : GEN_213;
  assign GEN_215 = 3'h7 == T_186_up_idx ? wmask_buffer_7 : GEN_214;
  assign T_3281 = {T_63,1'h0};
  assign T_3282 = {T_65,T_67};
  assign T_3283 = {T_3282,T_3281};
  assign T_3285 = {T_67,T_63};
  assign T_3286 = {T_3285,1'h0};
  assign T_3288 = {GEN_11,1'h0};
  assign T_3300 = T_2111 ? 6'h2 : {{5'd0}, 1'h0};
  assign T_3302 = T_2113 ? 6'h0 : T_3300;
  assign T_3304 = T_2109 ? T_3283 : {{6'd0}, T_3302};
  assign T_3306 = T_2119 ? {{3'd0}, T_3288} : T_3304;
  assign T_3308 = T_2115 ? {{3'd0}, T_3288} : T_3306;
  assign T_3310 = T_2121 ? {{3'd0}, T_3286} : T_3308;
  assign T_3312 = T_2117 ? T_3283 : T_3310;
  assign T_3341_addr_block = T_57;
  assign T_3341_client_xact_id = {{2'd0}, 1'h0};
  assign T_3341_addr_beat = T_186_up_idx;
  assign T_3341_is_builtin_type = 1'h1;
  assign T_3341_a_type = T_99_a_type;
  assign T_3341_union = T_3312;
  assign T_3341_data = GEN_12;
  assign GEN_12 = GEN_222;
  assign GEN_216 = GEN_444 == T_186_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_217 = GEN_465 == T_186_up_idx ? data_buffer_2 : GEN_216;
  assign GEN_218 = GEN_466 == T_186_up_idx ? data_buffer_3 : GEN_217;
  assign GEN_219 = 3'h4 == T_186_up_idx ? data_buffer_4 : GEN_218;
  assign GEN_220 = 3'h5 == T_186_up_idx ? data_buffer_5 : GEN_219;
  assign GEN_221 = 3'h6 == T_186_up_idx ? data_buffer_6 : GEN_220;
  assign GEN_222 = 3'h7 == T_186_up_idx ? data_buffer_7 : GEN_221;
  assign T_3369_addr_block = T_3074 ? T_3216_addr_block : T_3341_addr_block;
  assign T_3369_client_xact_id = T_3074 ? T_3216_client_xact_id : T_3341_client_xact_id;
  assign T_3369_addr_beat = T_3074 ? T_3216_addr_beat : T_3341_addr_beat;
  assign T_3369_is_builtin_type = T_3074 ? T_3216_is_builtin_type : T_3341_is_builtin_type;
  assign T_3369_a_type = T_3074 ? T_3216_a_type : T_3341_a_type;
  assign T_3369_union = T_3074 ? T_3216_union : T_3341_union;
  assign T_3369_data = T_3074 ? T_3216_data : T_3341_data;
  assign T_3398 = T_3162 & T_186_up_done;
  assign GEN_223 = T_3398 ? 4'h7 : GEN_55;
  assign T_3408_0 = 3'h5;
  assign T_3408_1 = 3'h4;
  assign GEN_527 = {{1'd0}, T_3408_0};
  assign T_3410 = GEN_527 == io_outer_grant_bits_g_type;
  assign GEN_528 = {{1'd0}, T_3408_1};
  assign T_3411 = GEN_528 == io_outer_grant_bits_g_type;
  assign T_3414 = T_3410 | T_3411;
  assign T_3420_0 = 1'h0;
  assign GEN_529 = {{3'd0}, T_3420_0};
  assign T_3422 = GEN_529 == io_outer_grant_bits_g_type;
  assign T_3425 = io_outer_grant_bits_is_builtin_type ? T_3414 : T_3422;
  assign T_3426 = T_2405 & T_3425;
  assign GEN_13 = GEN_230;
  assign GEN_224 = GEN_444 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_225 = GEN_465 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_224;
  assign GEN_226 = GEN_466 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_225;
  assign GEN_227 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_226;
  assign GEN_228 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_227;
  assign GEN_229 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_228;
  assign GEN_230 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_229;
  assign T_3427 = GEN_13[0];
  assign GEN_14 = GEN_230;
  assign T_3428 = GEN_14[1];
  assign GEN_15 = GEN_230;
  assign T_3429 = GEN_15[2];
  assign GEN_16 = GEN_230;
  assign T_3430 = GEN_16[3];
  assign GEN_17 = GEN_230;
  assign T_3431 = GEN_17[4];
  assign GEN_18 = GEN_230;
  assign T_3432 = GEN_18[5];
  assign GEN_19 = GEN_230;
  assign T_3433 = GEN_19[6];
  assign GEN_20 = GEN_230;
  assign T_3434 = GEN_20[7];
  assign GEN_554 = {{7'd0}, T_3427};
  assign T_3436 = 8'h0 - GEN_554;
  assign T_3437 = T_3436[7:0];
  assign GEN_555 = {{7'd0}, T_3428};
  assign T_3439 = 8'h0 - GEN_555;
  assign T_3440 = T_3439[7:0];
  assign GEN_556 = {{7'd0}, T_3429};
  assign T_3442 = 8'h0 - GEN_556;
  assign T_3443 = T_3442[7:0];
  assign GEN_557 = {{7'd0}, T_3430};
  assign T_3445 = 8'h0 - GEN_557;
  assign T_3446 = T_3445[7:0];
  assign GEN_558 = {{7'd0}, T_3431};
  assign T_3448 = 8'h0 - GEN_558;
  assign T_3449 = T_3448[7:0];
  assign GEN_559 = {{7'd0}, T_3432};
  assign T_3451 = 8'h0 - GEN_559;
  assign T_3452 = T_3451[7:0];
  assign GEN_560 = {{7'd0}, T_3433};
  assign T_3454 = 8'h0 - GEN_560;
  assign T_3455 = T_3454[7:0];
  assign GEN_561 = {{7'd0}, T_3434};
  assign T_3457 = 8'h0 - GEN_561;
  assign T_3458 = T_3457[7:0];
  assign T_3464_0 = T_3437;
  assign T_3464_1 = T_3440;
  assign T_3464_2 = T_3443;
  assign T_3464_3 = T_3446;
  assign T_3464_4 = T_3449;
  assign T_3464_5 = T_3452;
  assign T_3464_6 = T_3455;
  assign T_3464_7 = T_3458;
  assign T_3466 = {T_3464_1,T_3464_0};
  assign T_3467 = {T_3464_3,T_3464_2};
  assign T_3468 = {T_3467,T_3466};
  assign T_3469 = {T_3464_5,T_3464_4};
  assign T_3470 = {T_3464_7,T_3464_6};
  assign T_3471 = {T_3470,T_3469};
  assign T_3472 = {T_3471,T_3468};
  assign T_3473 = ~ T_3472;
  assign T_3474 = T_3473 & io_outer_grant_bits_data;
  assign GEN_21 = GEN_286;
  assign GEN_280 = GEN_444 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_281 = GEN_465 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_280;
  assign GEN_282 = GEN_466 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_281;
  assign GEN_283 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_282;
  assign GEN_284 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_283;
  assign GEN_285 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_284;
  assign GEN_286 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_285;
  assign T_3475 = T_3472 & GEN_21;
  assign T_3476 = T_3474 | T_3475;
  assign GEN_22 = T_3476;
  assign GEN_287 = GEN_433 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_177;
  assign GEN_288 = GEN_444 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_178;
  assign GEN_289 = GEN_465 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_179;
  assign GEN_290 = GEN_466 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_180;
  assign GEN_291 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_181;
  assign GEN_292 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_182;
  assign GEN_293 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_183;
  assign GEN_294 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_184;
  assign GEN_313 = T_3426 ? GEN_287 : GEN_177;
  assign GEN_314 = T_3426 ? GEN_288 : GEN_178;
  assign GEN_315 = T_3426 ? GEN_289 : GEN_179;
  assign GEN_316 = T_3426 ? GEN_290 : GEN_180;
  assign GEN_317 = T_3426 ? GEN_291 : GEN_181;
  assign GEN_318 = T_3426 ? GEN_292 : GEN_182;
  assign GEN_319 = T_3426 ? GEN_293 : GEN_183;
  assign GEN_320 = T_3426 ? GEN_294 : GEN_184;
  assign T_3477 = T_221 | T_186_pending;
  assign T_3478 = T_3477 | T_210_pending;
  assign T_3489 = T_2325 == 1'h0;
  assign T_3491 = T_2321 & T_3489;
  assign T_3499_0 = 3'h5;
  assign GEN_570 = {{1'd0}, T_3499_0};
  assign T_3501 = GEN_570 == io_inner_grant_bits_g_type;
  assign T_3509_0 = 2'h0;
  assign T_3509_1 = 2'h1;
  assign GEN_571 = {{2'd0}, T_3509_0};
  assign T_3511 = GEN_571 == io_inner_grant_bits_g_type;
  assign GEN_572 = {{2'd0}, T_3509_1};
  assign T_3512 = GEN_572 == io_inner_grant_bits_g_type;
  assign T_3515 = T_3511 | T_3512;
  assign T_3516 = io_inner_grant_bits_is_builtin_type ? T_3501 : T_3515;
  assign T_3518 = T_3491 & T_3516;
  assign T_3522 = T_3520 == 3'h7;
  assign T_3524 = T_3520 + GEN_444;
  assign T_3525 = T_3524[2:0];
  assign GEN_321 = T_3518 ? T_3525 : T_3520;
  assign T_3526 = T_3518 & T_3522;
  assign T_3527 = T_3516 ? T_3520 : {{2'd0}, 1'h0};
  assign T_3528 = T_3516 ? T_3526 : T_3491;
  assign T_3529 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3547 = T_3529 == 1'h0;
  assign T_3548 = T_3528 & T_3547;
  assign T_3550 = T_3545 + 1'h1;
  assign T_3551 = T_3550[0:0];
  assign GEN_323 = T_3548 ? T_3551 : T_3545;
  assign T_3553 = T_3528 == 1'h0;
  assign T_3554 = T_3529 & T_3553;
  assign T_3556 = T_3545 - 1'h1;
  assign T_3557 = T_3556[0:0];
  assign GEN_324 = T_3554 ? T_3557 : GEN_323;
  assign T_3559 = T_3545 > 1'h0;
  assign T_3564 = T_1885 == 1'h0;
  assign T_3573_0 = 3'h5;
  assign T_3573_1 = 3'h4;
  assign GEN_575 = {{1'd0}, T_3573_0};
  assign T_3575 = GEN_575 == io_inner_grant_bits_g_type;
  assign GEN_576 = {{1'd0}, T_3573_1};
  assign T_3576 = GEN_576 == io_inner_grant_bits_g_type;
  assign T_3579 = T_3575 | T_3576;
  assign T_3585_0 = 2'h0;
  assign T_3585_1 = 2'h1;
  assign GEN_577 = {{2'd0}, T_3585_0};
  assign T_3587 = GEN_577 == io_inner_grant_bits_g_type;
  assign GEN_578 = {{2'd0}, T_3585_1};
  assign T_3588 = GEN_578 == io_inner_grant_bits_g_type;
  assign T_3591 = T_3587 | T_3588;
  assign T_3592 = io_inner_grant_bits_is_builtin_type ? T_3579 : T_3591;
  assign T_3593 = T_2321 & T_3592;
  assign GEN_579 = {{7'd0}, T_3593};
  assign T_3595 = 8'h0 - GEN_579;
  assign T_3596 = T_3595[7:0];
  assign T_3597 = ~ T_3596;
  assign T_3599 = GEN_437 << io_inner_grant_bits_addr_beat;
  assign T_3600 = ~ T_3599;
  assign T_3601 = T_3597 | T_3600;
  assign T_3602 = T_177 & T_3601;
  assign T_3610_0 = 3'h0;
  assign T_3610_1 = 3'h1;
  assign T_3610_2 = 3'h2;
  assign T_3612 = T_3610_0 == io_inner_release_bits_r_type;
  assign T_3613 = T_3610_1 == io_inner_release_bits_r_type;
  assign T_3614 = T_3610_2 == io_inner_release_bits_r_type;
  assign T_3617 = T_3612 | T_3613;
  assign T_3618 = T_3617 | T_3614;
  assign T_3619 = T_2228 & T_3618;
  assign GEN_581 = {{7'd0}, T_3619};
  assign T_3622 = 8'h0 - GEN_581;
  assign T_3623 = T_3622[7:0];
  assign T_3626 = T_3623 & T_2476;
  assign T_3627 = T_3602 | T_3626;
  assign T_3637_0 = 3'h5;
  assign T_3637_1 = 3'h4;
  assign GEN_583 = {{1'd0}, T_3637_0};
  assign T_3639 = GEN_583 == io_outer_grant_bits_g_type;
  assign GEN_584 = {{1'd0}, T_3637_1};
  assign T_3640 = GEN_584 == io_outer_grant_bits_g_type;
  assign T_3643 = T_3639 | T_3640;
  assign T_3649_0 = 1'h0;
  assign GEN_585 = {{3'd0}, T_3649_0};
  assign T_3651 = GEN_585 == io_outer_grant_bits_g_type;
  assign T_3654 = io_outer_grant_bits_is_builtin_type ? T_3643 : T_3651;
  assign T_3655 = T_2405 & T_3654;
  assign GEN_586 = {{7'd0}, T_3655};
  assign T_3658 = 8'h0 - GEN_586;
  assign T_3659 = T_3658[7:0];
  assign T_3661 = GEN_437 << io_outer_grant_bits_addr_beat;
  assign T_3662 = T_3659 & T_3661;
  assign T_3663 = T_3627 | T_3662;
  assign T_3664 = T_3663 | GEN_432;
  assign GEN_335 = T_3564 ? T_3664 : GEN_43;
  assign T_3666 = T_55 == 4'h1;
  assign T_3667 = T_1733 | T_3666;
  assign T_3670 = T_3667 | T_2075;
  assign T_3672 = T_3670 == 1'h0;
  assign T_3689 = 3'h6 == Queue_12_1_io_deq_bits_a_type;
  assign T_3690 = T_3689 ? 3'h1 : 3'h3;
  assign T_3691 = 3'h5 == Queue_12_1_io_deq_bits_a_type;
  assign T_3692 = T_3691 ? 3'h1 : T_3690;
  assign T_3693 = 3'h4 == Queue_12_1_io_deq_bits_a_type;
  assign T_3694 = T_3693 ? 3'h4 : T_3692;
  assign T_3695 = 3'h3 == Queue_12_1_io_deq_bits_a_type;
  assign T_3696 = T_3695 ? 3'h3 : T_3694;
  assign T_3697 = 3'h2 == Queue_12_1_io_deq_bits_a_type;
  assign T_3698 = T_3697 ? 3'h3 : T_3696;
  assign T_3699 = 3'h1 == Queue_12_1_io_deq_bits_a_type;
  assign T_3700 = T_3699 ? 3'h5 : T_3698;
  assign T_3701 = 3'h0 == Queue_12_1_io_deq_bits_a_type;
  assign T_3702 = T_3701 ? 3'h4 : T_3700;
  assign T_3703 = Queue_12_1_io_deq_bits_a_type == GEN_433;
  assign T_3708 = T_3703 ? 2'h0 : 2'h1;
  assign T_3709 = Queue_12_1_io_deq_bits_is_builtin_type ? T_3702 : {{1'd0}, T_3708};
  assign T_3741_addr_beat = Queue_12_1_io_deq_bits_addr_beat;
  assign T_3741_client_xact_id = Queue_12_1_io_deq_bits_client_xact_id;
  assign T_3741_manager_xact_id = {{1'd0}, 2'h2};
  assign T_3741_is_builtin_type = Queue_12_1_io_deq_bits_is_builtin_type;
  assign T_3741_g_type = {{1'd0}, T_3709};
  assign T_3741_data = GEN_23;
  assign T_3741_client_id = Queue_12_1_io_deq_bits_client_id;
  assign GEN_23 = GEN_342;
  assign GEN_336 = GEN_444 == T_155 ? data_buffer_1 : data_buffer_0;
  assign GEN_337 = GEN_465 == T_155 ? data_buffer_2 : GEN_336;
  assign GEN_338 = GEN_466 == T_155 ? data_buffer_3 : GEN_337;
  assign GEN_339 = 3'h4 == T_155 ? data_buffer_4 : GEN_338;
  assign GEN_340 = 3'h5 == T_155 ? data_buffer_5 : GEN_339;
  assign GEN_341 = 3'h6 == T_155 ? data_buffer_6 : GEN_340;
  assign GEN_342 = 3'h7 == T_155 ? data_buffer_7 : GEN_341;
  assign T_3780_0 = 3'h5;
  assign GEN_594 = {{1'd0}, T_3780_0};
  assign T_3782 = GEN_594 == io_inner_grant_bits_g_type;
  assign T_3790_0 = 2'h0;
  assign T_3790_1 = 2'h1;
  assign GEN_595 = {{2'd0}, T_3790_0};
  assign T_3792 = GEN_595 == io_inner_grant_bits_g_type;
  assign GEN_596 = {{2'd0}, T_3790_1};
  assign T_3793 = GEN_596 == io_inner_grant_bits_g_type;
  assign T_3796 = T_3792 | T_3793;
  assign T_3797 = io_inner_grant_bits_is_builtin_type ? T_3782 : T_3796;
  assign T_3799 = T_2321 & T_3797;
  assign T_3803 = T_3801 == 3'h7;
  assign T_3805 = T_3801 + GEN_444;
  assign T_3806 = T_3805[2:0];
  assign GEN_343 = T_3799 ? T_3806 : T_3801;
  assign T_3807 = T_3799 & T_3803;
  assign T_3808 = T_3797 ? T_3801 : Queue_12_1_io_deq_bits_addr_beat;
  assign T_3809 = T_3797 ? T_3807 : T_2321;
  assign T_3814 = T_2977 & T_153;
  assign T_3816 = T_3478 == 1'h0;
  assign T_3824_0 = 3'h5;
  assign T_3824_1 = 3'h4;
  assign GEN_598 = {{1'd0}, T_3824_0};
  assign T_3826 = GEN_598 == io_inner_grant_bits_g_type;
  assign GEN_599 = {{1'd0}, T_3824_1};
  assign T_3827 = GEN_599 == io_inner_grant_bits_g_type;
  assign T_3830 = T_3826 | T_3827;
  assign T_3836_0 = 2'h0;
  assign T_3836_1 = 2'h1;
  assign GEN_600 = {{2'd0}, T_3836_0};
  assign T_3838 = GEN_600 == io_inner_grant_bits_g_type;
  assign GEN_601 = {{2'd0}, T_3836_1};
  assign T_3839 = GEN_601 == io_inner_grant_bits_g_type;
  assign T_3842 = T_3838 | T_3839;
  assign T_3843 = io_inner_grant_bits_is_builtin_type ? T_3830 : T_3842;
  assign T_3844 = T_177 >> T_155;
  assign T_3845 = T_3844[0];
  assign T_3846 = T_3843 ? T_3845 : T_3672;
  assign T_3847 = T_3816 & T_3846;
  assign GEN_348 = T_3814 ? T_3847 : T_2537;
  assign GEN_349 = T_2414 ? T_157 : 1'h0;
  assign GEN_350 = T_2414 ? T_155 : T_2639_addr_beat;
  assign GEN_351 = T_2414 ? T_3741_client_xact_id : T_2639_client_xact_id;
  assign GEN_352 = T_2414 ? T_3741_manager_xact_id : T_2639_manager_xact_id;
  assign GEN_353 = T_2414 ? T_3741_is_builtin_type : T_2639_is_builtin_type;
  assign GEN_354 = T_2414 ? T_3741_g_type : T_2639_g_type;
  assign GEN_355 = T_2414 ? T_3741_data : T_2639_data;
  assign GEN_356 = T_2414 ? T_3741_client_id : T_2639_client_id;
  assign GEN_361 = T_2414 ? GEN_348 : T_2537;
  assign T_3854 = ~ io_incoherent_0;
  assign GEN_362 = T_1885 ? {{1'd0}, T_3854} : T_2207;
  assign T_3869_0 = 3'h3;
  assign T_3871 = T_3869_0 == T_99_a_type;
  assign T_3874 = T_99_is_builtin_type & T_3871;
  assign T_3875 = T_1887 & T_3874;
  assign T_3876 = T_3875 & T_153;
  assign T_3879 = T_3876 & T_1905;
  assign T_3881 = T_3879 & io_inner_acquire_valid;
  assign T_3882 = T_1885 | T_3881;
  assign T_3892_0 = 3'h2;
  assign T_3892_1 = 3'h3;
  assign T_3892_2 = 3'h4;
  assign T_3894 = T_3892_0 == io_inner_acquire_bits_a_type;
  assign T_3895 = T_3892_1 == io_inner_acquire_bits_a_type;
  assign T_3896 = T_3892_2 == io_inner_acquire_bits_a_type;
  assign T_3899 = T_3894 | T_3895;
  assign T_3900 = T_3899 | T_3896;
  assign T_3901 = io_inner_acquire_bits_is_builtin_type & T_3900;
  assign T_3902 = T_1734 & T_3901;
  assign T_3903 = T_3902 & T_3882;
  assign T_3905 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3906 = io_inner_acquire_bits_is_builtin_type & T_3905;
  assign T_3910 = 8'h0 - GEN_437;
  assign T_3911 = T_3910[7:0];
  assign T_3917_0 = T_3911;
  assign T_3925 = T_2034 | T_2031;
  assign T_3926 = io_inner_acquire_bits_union[8:1];
  assign T_3928 = T_3925 ? T_3926 : {{7'd0}, 1'h0};
  assign T_3929 = T_3906 ? T_3917_0 : T_3928;
  assign T_3930 = T_3929[0];
  assign T_3931 = T_3929[1];
  assign T_3932 = T_3929[2];
  assign T_3933 = T_3929[3];
  assign T_3934 = T_3929[4];
  assign T_3935 = T_3929[5];
  assign T_3936 = T_3929[6];
  assign T_3937 = T_3929[7];
  assign GEN_603 = {{7'd0}, T_3930};
  assign T_3939 = 8'h0 - GEN_603;
  assign T_3940 = T_3939[7:0];
  assign GEN_604 = {{7'd0}, T_3931};
  assign T_3942 = 8'h0 - GEN_604;
  assign T_3943 = T_3942[7:0];
  assign GEN_605 = {{7'd0}, T_3932};
  assign T_3945 = 8'h0 - GEN_605;
  assign T_3946 = T_3945[7:0];
  assign GEN_606 = {{7'd0}, T_3933};
  assign T_3948 = 8'h0 - GEN_606;
  assign T_3949 = T_3948[7:0];
  assign GEN_607 = {{7'd0}, T_3934};
  assign T_3951 = 8'h0 - GEN_607;
  assign T_3952 = T_3951[7:0];
  assign GEN_608 = {{7'd0}, T_3935};
  assign T_3954 = 8'h0 - GEN_608;
  assign T_3955 = T_3954[7:0];
  assign GEN_609 = {{7'd0}, T_3936};
  assign T_3957 = 8'h0 - GEN_609;
  assign T_3958 = T_3957[7:0];
  assign GEN_610 = {{7'd0}, T_3937};
  assign T_3960 = 8'h0 - GEN_610;
  assign T_3961 = T_3960[7:0];
  assign T_3967_0 = T_3940;
  assign T_3967_1 = T_3943;
  assign T_3967_2 = T_3946;
  assign T_3967_3 = T_3949;
  assign T_3967_4 = T_3952;
  assign T_3967_5 = T_3955;
  assign T_3967_6 = T_3958;
  assign T_3967_7 = T_3961;
  assign T_3969 = {T_3967_1,T_3967_0};
  assign T_3970 = {T_3967_3,T_3967_2};
  assign T_3971 = {T_3970,T_3969};
  assign T_3972 = {T_3967_5,T_3967_4};
  assign T_3973 = {T_3967_7,T_3967_6};
  assign T_3974 = {T_3973,T_3972};
  assign T_3975 = {T_3974,T_3971};
  assign T_3976 = ~ T_3975;
  assign GEN_24 = GEN_369;
  assign GEN_363 = GEN_444 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_364 = GEN_465 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_363;
  assign GEN_365 = GEN_466 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_364;
  assign GEN_366 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_365;
  assign GEN_367 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_366;
  assign GEN_368 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_367;
  assign GEN_369 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_368;
  assign T_3977 = T_3976 & GEN_24;
  assign T_3978 = T_3975 & io_inner_acquire_bits_data;
  assign T_3979 = T_3977 | T_3978;
  assign GEN_25 = T_3979;
  assign GEN_370 = GEN_433 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_313;
  assign GEN_371 = GEN_444 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_314;
  assign GEN_372 = GEN_465 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_315;
  assign GEN_373 = GEN_466 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_316;
  assign GEN_374 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_317;
  assign GEN_375 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_318;
  assign GEN_376 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_319;
  assign GEN_377 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_320;
  assign T_3993_0 = T_3911;
  assign T_4005 = T_3906 ? T_3993_0 : T_3928;
  assign GEN_26 = GEN_384;
  assign GEN_378 = GEN_444 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_379 = GEN_465 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_378;
  assign GEN_380 = GEN_466 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_379;
  assign GEN_381 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_380;
  assign GEN_382 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_381;
  assign GEN_383 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_382;
  assign GEN_384 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_383;
  assign T_4006 = T_4005 | GEN_26;
  assign GEN_27 = T_4006;
  assign GEN_385 = GEN_433 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_0;
  assign GEN_386 = GEN_444 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_1;
  assign GEN_387 = GEN_465 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_2;
  assign GEN_388 = GEN_466 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_3;
  assign GEN_389 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_4;
  assign GEN_390 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_5;
  assign GEN_391 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_6;
  assign GEN_392 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_7;
  assign GEN_404 = T_3903 ? GEN_370 : GEN_313;
  assign GEN_405 = T_3903 ? GEN_371 : GEN_314;
  assign GEN_406 = T_3903 ? GEN_372 : GEN_315;
  assign GEN_407 = T_3903 ? GEN_373 : GEN_316;
  assign GEN_408 = T_3903 ? GEN_374 : GEN_317;
  assign GEN_409 = T_3903 ? GEN_375 : GEN_318;
  assign GEN_410 = T_3903 ? GEN_376 : GEN_319;
  assign GEN_411 = T_3903 ? GEN_377 : GEN_320;
  assign GEN_415 = T_3903 ? GEN_385 : wmask_buffer_0;
  assign GEN_416 = T_3903 ? GEN_386 : wmask_buffer_1;
  assign GEN_417 = T_3903 ? GEN_387 : wmask_buffer_2;
  assign GEN_418 = T_3903 ? GEN_388 : wmask_buffer_3;
  assign GEN_419 = T_3903 ? GEN_389 : wmask_buffer_4;
  assign GEN_420 = T_3903 ? GEN_390 : wmask_buffer_5;
  assign GEN_421 = T_3903 ? GEN_391 : wmask_buffer_6;
  assign GEN_422 = T_3903 ? GEN_392 : wmask_buffer_7;
  assign T_4009 = T_2075 | T_2533;
  assign T_4010 = T_4009 | T_144_pending;
  assign T_4011 = T_4010 | T_221;
  assign T_4012 = T_4011 | T_210_pending;
  assign T_4013 = T_4012 | T_186_pending;
  assign T_4014 = T_4013 | T_153;
  assign T_4015 = T_4014 | T_166_pending;
  assign T_4017 = T_4015 == 1'h0;
  assign T_4019 = T_2977 & T_44;
  assign GEN_423 = T_4019 ? 4'h0 : GEN_223;
  assign GEN_424 = T_4019 ? {{7'd0}, 1'h0} : GEN_415;
  assign GEN_425 = T_4019 ? {{7'd0}, 1'h0} : GEN_416;
  assign GEN_426 = T_4019 ? {{7'd0}, 1'h0} : GEN_417;
  assign GEN_427 = T_4019 ? {{7'd0}, 1'h0} : GEN_418;
  assign GEN_428 = T_4019 ? {{7'd0}, 1'h0} : GEN_419;
  assign GEN_429 = T_4019 ? {{7'd0}, 1'h0} : GEN_420;
  assign GEN_430 = T_4019 ? {{7'd0}, 1'h0} : GEN_421;
  assign GEN_431 = T_4019 ? {{7'd0}, 1'h0} : GEN_422;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_30 = {1{$random}};
  T_55 = GEN_30[3:0];
  GEN_31 = {1{$random}};
  T_57 = GEN_31[25:0];
  GEN_39 = {1{$random}};
  T_59 = GEN_39[0:0];
  GEN_40 = {1{$random}};
  T_61 = GEN_40[4:0];
  GEN_41 = {1{$random}};
  T_63 = GEN_41[4:0];
  GEN_45 = {1{$random}};
  T_65 = GEN_45[2:0];
  GEN_59 = {1{$random}};
  T_67 = GEN_59[2:0];
  GEN_60 = {1{$random}};
  T_129 = GEN_60[2:0];
  GEN_61 = {1{$random}};
  T_131 = GEN_61[0:0];
  GEN_62 = {1{$random}};
  T_133 = GEN_62[1:0];
  GEN_63 = {1{$random}};
  T_135 = GEN_63[7:0];
  GEN_64 = {1{$random}};
  T_175 = GEN_64[7:0];
  GEN_66 = {1{$random}};
  T_177 = GEN_66[7:0];
  GEN_67 = {1{$random}};
  T_195 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  T_199 = GEN_68[0:0];
  GEN_70 = {1{$random}};
  T_201 = GEN_70[7:0];
  GEN_71 = {2{$random}};
  data_buffer_0 = GEN_71[63:0];
  GEN_72 = {2{$random}};
  data_buffer_1 = GEN_72[63:0];
  GEN_73 = {2{$random}};
  data_buffer_2 = GEN_73[63:0];
  GEN_74 = {2{$random}};
  data_buffer_3 = GEN_74[63:0];
  GEN_78 = {2{$random}};
  data_buffer_4 = GEN_78[63:0];
  GEN_79 = {2{$random}};
  data_buffer_5 = GEN_79[63:0];
  GEN_80 = {2{$random}};
  data_buffer_6 = GEN_80[63:0];
  GEN_81 = {2{$random}};
  data_buffer_7 = GEN_81[63:0];
  GEN_82 = {1{$random}};
  wmask_buffer_0 = GEN_82[7:0];
  GEN_83 = {1{$random}};
  wmask_buffer_1 = GEN_83[7:0];
  GEN_85 = {1{$random}};
  wmask_buffer_2 = GEN_85[7:0];
  GEN_86 = {1{$random}};
  wmask_buffer_3 = GEN_86[7:0];
  GEN_87 = {1{$random}};
  wmask_buffer_4 = GEN_87[7:0];
  GEN_95 = {1{$random}};
  wmask_buffer_5 = GEN_95[7:0];
  GEN_96 = {1{$random}};
  wmask_buffer_6 = GEN_96[7:0];
  GEN_97 = {1{$random}};
  wmask_buffer_7 = GEN_97[7:0];
  GEN_98 = {1{$random}};
  T_2219 = GEN_98[2:0];
  GEN_99 = {1{$random}};
  T_2252 = GEN_99[2:0];
  GEN_100 = {1{$random}};
  T_2262 = GEN_100[0:0];
  GEN_101 = {1{$random}};
  T_2312 = GEN_101[2:0];
  GEN_102 = {1{$random}};
  T_2356 = GEN_102[2:0];
  GEN_103 = {1{$random}};
  T_2366 = GEN_103[0:0];
  GEN_104 = {1{$random}};
  T_2912 = GEN_104[2:0];
  GEN_105 = {1{$random}};
  T_2952 = GEN_105[2:0];
  GEN_106 = {1{$random}};
  T_2962 = GEN_106[0:0];
  GEN_107 = {1{$random}};
  T_3095 = GEN_107[2:0];
  GEN_108 = {1{$random}};
  T_3137 = GEN_108[2:0];
  GEN_109 = {1{$random}};
  T_3147 = GEN_109[0:0];
  GEN_110 = {1{$random}};
  T_3520 = GEN_110[2:0];
  GEN_111 = {1{$random}};
  T_3535 = GEN_111[2:0];
  GEN_112 = {1{$random}};
  T_3545 = GEN_112[0:0];
  GEN_113 = {1{$random}};
  T_3801 = GEN_113[2:0];
  GEN_114 = {1{$random}};
  GEN_28 = GEN_114[0:0];
  GEN_115 = {1{$random}};
  GEN_29 = GEN_115[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_55 <= 4'h0;
    end else begin
      if(T_4019) begin
        T_55 <= 4'h0;
      end else begin
        if(T_3398) begin
          T_55 <= 4'h7;
        end else begin
          if(T_2383) begin
            T_55 <= 4'h7;
          end else begin
            if(T_2283) begin
              if(T_2183) begin
                T_55 <= 4'h6;
              end else begin
                T_55 <= 4'h7;
              end
            end else begin
              if(T_1885) begin
                T_55 <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_57 <= 26'h0;
    end else begin
      if(T_2383) begin
        T_57 <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1885) begin
          T_57 <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_59 <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_61 <= T_2028;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        if(T_2035) begin
          T_63 <= 5'h1;
        end else begin
          T_63 <= T_2036;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_65 <= T_2038;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_67 <= T_2039;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_129 <= io_inner_release_bits_r_type;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_131 <= io_inner_release_bits_client_id;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_133 <= io_inner_release_bits_client_xact_id;
        end
      end
    end
    if(reset) begin
      T_135 <= 8'h0;
    end else begin
      if(T_2228) begin
        if(T_2489) begin
          T_135 <= T_2514;
        end else begin
          if(T_2438) begin
            if(T_2453) begin
              T_135 <= T_2478;
            end else begin
              T_135 <= {{7'd0}, 1'h0};
            end
          end
        end
      end
    end
    if(reset) begin
      T_175 <= 8'h0;
    end else begin
      if(T_1885) begin
        if(T_2034) begin
          T_175 <= T_2070;
        end else begin
          T_175 <= {{7'd0}, 1'h0};
        end
      end else begin
        if(T_1962) begin
          T_175 <= T_2020;
        end
      end
    end
    if(reset) begin
      T_177 <= 8'h0;
    end else begin
      if(T_3564) begin
        T_177 <= T_3664;
      end else begin
        if(T_1885) begin
          T_177 <= {{7'd0}, 1'h0};
        end
      end
    end
    if(1'h0) begin
    end else begin
      T_195 <= GEN_362[0];
    end
    if(reset) begin
      T_199 <= 1'h0;
    end else begin
      if(T_2833) begin
        T_199 <= 1'h0;
      end
    end
    if(reset) begin
      T_201 <= 8'h0;
    end else begin
      if(T_2832) begin
        T_201 <= T_2883;
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1817_0;
    end else begin
      if(T_3903) begin
        if(GEN_433 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_433 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_433 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_433 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_433 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_433 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_433 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1817_1;
    end else begin
      if(T_3903) begin
        if(GEN_444 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_444 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_444 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_444 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_444 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_444 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_444 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1817_2;
    end else begin
      if(T_3903) begin
        if(GEN_465 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_465 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_465 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_465 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_465 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_465 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_465 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1817_3;
    end else begin
      if(T_3903) begin
        if(GEN_466 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_466 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_466 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_466 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_466 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_466 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_466 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1817_4;
    end else begin
      if(T_3903) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1817_5;
    end else begin
      if(T_3903) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1817_6;
    end else begin
      if(T_3903) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1817_7;
    end else begin
      if(T_3903) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1835_0;
    end else begin
      if(T_4019) begin
        wmask_buffer_0 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_433 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1835_1;
    end else begin
      if(T_4019) begin
        wmask_buffer_1 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_444 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1835_2;
    end else begin
      if(T_4019) begin
        wmask_buffer_2 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_465 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1835_3;
    end else begin
      if(T_4019) begin
        wmask_buffer_3 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_466 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1835_4;
    end else begin
      if(T_4019) begin
        wmask_buffer_4 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1835_5;
    end else begin
      if(T_4019) begin
        wmask_buffer_5 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1835_6;
    end else begin
      if(T_4019) begin
        wmask_buffer_6 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1835_7;
    end else begin
      if(T_4019) begin
        wmask_buffer_7 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      T_2219 <= 3'h0;
    end
    if(reset) begin
      T_2252 <= 3'h0;
    end else begin
      if(T_2250) begin
        T_2252 <= T_2257;
      end
    end
    if(reset) begin
      T_2262 <= 1'h0;
    end else begin
      if(T_2271) begin
        T_2262 <= T_2274;
      end else begin
        if(T_2265) begin
          T_2262 <= T_2268;
        end
      end
    end
    if(reset) begin
      T_2312 <= 3'h0;
    end else begin
      if(T_2310) begin
        T_2312 <= T_2317;
      end
    end
    if(reset) begin
      T_2356 <= 3'h0;
    end else begin
      if(T_2354) begin
        T_2356 <= T_2361;
      end
    end
    if(reset) begin
      T_2366 <= 1'h0;
    end else begin
      if(T_2375) begin
        T_2366 <= T_2378;
      end else begin
        if(T_2369) begin
          T_2366 <= T_2372;
        end
      end
    end
    if(reset) begin
      T_2912 <= 3'h0;
    end else begin
      if(T_2910) begin
        T_2912 <= T_2917;
      end
    end
    if(reset) begin
      T_2952 <= 3'h0;
    end else begin
      if(T_2950) begin
        T_2952 <= T_2957;
      end
    end
    if(reset) begin
      T_2962 <= 1'h0;
    end else begin
      if(T_2971) begin
        T_2962 <= T_2974;
      end else begin
        if(T_2965) begin
          T_2962 <= T_2968;
        end
      end
    end
    if(reset) begin
      T_3095 <= 3'h0;
    end else begin
      if(T_3093) begin
        T_3095 <= T_3100;
      end
    end
    if(reset) begin
      T_3137 <= 3'h0;
    end else begin
      if(T_3135) begin
        T_3137 <= T_3142;
      end
    end
    if(reset) begin
      T_3147 <= 1'h0;
    end else begin
      if(T_3156) begin
        T_3147 <= T_3159;
      end else begin
        if(T_3150) begin
          T_3147 <= T_3153;
        end
      end
    end
    if(reset) begin
      T_3520 <= 3'h0;
    end else begin
      if(T_3518) begin
        T_3520 <= T_3525;
      end
    end
    if(reset) begin
      T_3535 <= 3'h0;
    end
    if(reset) begin
      T_3545 <= 1'h0;
    end else begin
      if(T_3554) begin
        T_3545 <= T_3557;
      end else begin
        if(T_3548) begin
          T_3545 <= T_3551;
        end
      end
    end
    if(reset) begin
      T_3801 <= 3'h0;
    end else begin
      if(T_3799) begin
        T_3801 <= T_3806;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1778) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:95 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1778) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1778) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1792) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:99 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1792) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1792) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1803) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1803) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1803) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BufferedBroadcastAcquireTracker_2(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should
);
  wire  T_44;
  reg [3:0] T_55;
  reg [31:0] GEN_30;
  reg [25:0] T_57;
  reg [31:0] GEN_31;
  reg  T_59;
  reg [31:0] GEN_39;
  reg [4:0] T_61;
  reg [31:0] GEN_40;
  reg [4:0] T_63;
  reg [31:0] GEN_41;
  reg [2:0] T_65;
  reg [31:0] GEN_45;
  reg [2:0] T_67;
  reg [31:0] GEN_59;
  wire [2:0] T_69;
  wire [1:0] T_99_client_xact_id;
  wire [2:0] T_99_addr_beat;
  wire  T_99_client_id;
  wire  T_99_is_builtin_type;
  wire [2:0] T_99_a_type;
  reg [2:0] T_129;
  reg [31:0] GEN_60;
  reg  T_131;
  reg [31:0] GEN_61;
  reg [1:0] T_133;
  reg [31:0] GEN_62;
  reg [7:0] T_135;
  reg [31:0] GEN_63;
  wire  T_144_pending;
  wire [2:0] T_144_up_idx;
  wire  T_144_up_done;
  wire [2:0] T_144_down_idx;
  wire  T_144_down_done;
  wire  T_153;
  wire [2:0] T_155;
  wire  T_157;
  wire  T_166_pending;
  wire [2:0] T_166_up_idx;
  wire  T_166_up_done;
  wire [2:0] T_166_down_idx;
  wire  T_166_down_done;
  reg [7:0] T_175;
  reg [31:0] GEN_64;
  reg [7:0] T_177;
  reg [31:0] GEN_66;
  wire  T_186_pending;
  wire [2:0] T_186_up_idx;
  wire  T_186_up_done;
  wire [2:0] T_186_down_idx;
  wire  T_186_down_done;
  reg  T_195;
  reg [31:0] GEN_67;
  reg  T_199;
  reg [31:0] GEN_68;
  reg [7:0] T_201;
  reg [31:0] GEN_70;
  wire  T_210_pending;
  wire [2:0] T_210_up_idx;
  wire  T_210_up_done;
  wire [2:0] T_210_down_idx;
  wire  T_210_down_done;
  wire [7:0] GEN_432;
  wire  T_219;
  wire  T_220;
  wire  T_221;
  wire  T_247_sharers;
  wire [1:0] T_299_state;
  wire  T_395_inner_sharers;
  wire [1:0] T_395_outer_state;
  wire  T_1733;
  wire  T_1734;
  wire  T_1735;
  wire  T_1736;
  wire [2:0] T_1745_0;
  wire  T_1747;
  wire  T_1750;
  wire  T_1751;
  wire [2:0] T_1760_0;
  wire  T_1762;
  wire  T_1765;
  wire  T_1767;
  wire [2:0] GEN_433;
  wire  T_1769;
  wire  T_1770;
  wire  T_1772;
  wire  T_1773;
  wire  T_1775;
  wire  T_1776;
  wire  T_1778;
  wire  T_1779;
  wire  T_1780;
  wire  T_1782;
  wire  T_1784;
  wire  T_1785;
  wire  T_1786;
  wire  T_1787;
  wire  T_1789;
  wire  T_1790;
  wire  T_1792;
  wire  T_1796;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [63:0] T_1817_0;
  wire [63:0] T_1817_1;
  wire [63:0] T_1817_2;
  wire [63:0] T_1817_3;
  wire [63:0] T_1817_4;
  wire [63:0] T_1817_5;
  wire [63:0] T_1817_6;
  wire [63:0] T_1817_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_71;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_72;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_73;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_74;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_78;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_79;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_80;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_81;
  wire [7:0] T_1835_0;
  wire [7:0] T_1835_1;
  wire [7:0] T_1835_2;
  wire [7:0] T_1835_3;
  wire [7:0] T_1835_4;
  wire [7:0] T_1835_5;
  wire [7:0] T_1835_6;
  wire [7:0] T_1835_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_82;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_83;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_85;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_86;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_87;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_95;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_96;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_97;
  wire  T_1841;
  wire  T_1842;
  wire  T_1844;
  wire  T_1845;
  wire  T_1847;
  wire  T_1848;
  wire  Queue_13_1_clk;
  wire  Queue_13_1_reset;
  wire  Queue_13_1_io_enq_ready;
  wire  Queue_13_1_io_enq_valid;
  wire [1:0] Queue_13_1_io_enq_bits_client_xact_id;
  wire [2:0] Queue_13_1_io_enq_bits_addr_beat;
  wire  Queue_13_1_io_enq_bits_client_id;
  wire  Queue_13_1_io_enq_bits_is_builtin_type;
  wire [2:0] Queue_13_1_io_enq_bits_a_type;
  wire  Queue_13_1_io_deq_ready;
  wire  Queue_13_1_io_deq_valid;
  wire [1:0] Queue_13_1_io_deq_bits_client_xact_id;
  wire [2:0] Queue_13_1_io_deq_bits_addr_beat;
  wire  Queue_13_1_io_deq_bits_client_id;
  wire  Queue_13_1_io_deq_bits_is_builtin_type;
  wire [2:0] Queue_13_1_io_deq_bits_a_type;
  wire [1:0] Queue_13_1_io_count;
  wire  T_1884;
  wire  T_1885;
  wire  T_1887;
  wire [2:0] T_1896_0;
  wire  T_1898;
  wire  T_1901;
  wire  T_1902;
  wire  T_1903;
  wire [7:0] T_1904;
  wire  T_1905;
  wire  T_1906;
  wire  T_1908;
  wire [2:0] T_1917_0;
  wire  T_1919;
  wire  T_1922;
  wire  T_1924;
  wire  T_1927;
  wire  T_1928;
  wire  T_1929;
  wire [1:0] T_1930_client_xact_id;
  wire [2:0] T_1930_addr_beat;
  wire  T_1930_client_id;
  wire  T_1930_is_builtin_type;
  wire [2:0] T_1930_a_type;
  wire [1:0] GEN_435;
  wire  T_1960;
  wire  T_1962;
  wire [2:0] T_1972_0;
  wire [2:0] T_1972_1;
  wire [2:0] T_1972_2;
  wire  T_1974;
  wire  T_1975;
  wire  T_1976;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire  T_1982;
  wire [7:0] GEN_436;
  wire [8:0] T_1984;
  wire [7:0] T_1985;
  wire [7:0] T_1986;
  wire [7:0] GEN_437;
  wire [7:0] T_1988;
  wire [7:0] T_1989;
  wire [7:0] T_1990;
  wire [7:0] T_1991;
  wire [2:0] T_2001_0;
  wire  T_2003;
  wire  T_2006;
  wire  T_2007;
  wire  T_2010;
  wire [7:0] T_2019;
  wire [7:0] T_2020;
  wire [7:0] GEN_32;
  wire [3:0] GEN_439;
  wire [4:0] T_2028;
  wire  T_2030;
  wire  T_2031;
  wire  T_2033;
  wire  T_2034;
  wire  T_2035;
  wire [4:0] T_2036;
  wire [4:0] T_2037;
  wire [2:0] T_2038;
  wire [2:0] T_2039;
  wire [2:0] T_2052_0;
  wire [2:0] T_2052_1;
  wire [2:0] T_2052_2;
  wire  T_2054;
  wire  T_2055;
  wire  T_2056;
  wire  T_2059;
  wire  T_2060;
  wire  T_2061;
  wire  T_2062;
  wire [7:0] GEN_440;
  wire [8:0] T_2064;
  wire [7:0] T_2065;
  wire [7:0] T_2066;
  wire [7:0] T_2070;
  wire [7:0] T_2072;
  wire [25:0] GEN_33;
  wire  GEN_34;
  wire [4:0] GEN_35;
  wire [4:0] GEN_36;
  wire [2:0] GEN_37;
  wire [2:0] GEN_38;
  wire [7:0] GEN_42;
  wire [7:0] GEN_43;
  wire [3:0] GEN_44;
  wire  T_2075;
  wire [2:0] T_2088_0;
  wire  T_2090;
  wire  T_2093;
  wire  T_2094;
  wire  T_2095;
  wire  T_2098;
  wire  T_2099;
  wire [7:0] T_2100;
  wire  skip_outer_acquire;
  wire  T_2109;
  wire [1:0] T_2110;
  wire  T_2111;
  wire [1:0] T_2112;
  wire  T_2113;
  wire [1:0] T_2114;
  wire  T_2115;
  wire [1:0] T_2116;
  wire  T_2117;
  wire [1:0] T_2118;
  wire  T_2119;
  wire [1:0] T_2120;
  wire  T_2121;
  wire [1:0] T_2122;
  wire [2:0] GEN_444;
  wire  T_2123;
  wire [1:0] T_2124;
  wire  T_2125;
  wire [1:0] T_2126;
  wire [1:0] T_2127;
  wire [25:0] T_2155_addr_block;
  wire [1:0] T_2155_p_type;
  wire  T_2155_client_id;
  wire  T_2183;
  wire [3:0] T_2184;
  wire  T_2193_pending;
  wire [2:0] T_2193_up_idx;
  wire  T_2193_up_done;
  wire [2:0] T_2193_down_idx;
  wire  T_2193_down_done;
  wire  T_2201;
  wire  T_2202;
  wire [1:0] GEN_446;
  wire [1:0] T_2204;
  wire [1:0] T_2205;
  wire [1:0] GEN_447;
  wire [1:0] T_2206;
  wire [1:0] GEN_448;
  wire [1:0] T_2207;
  wire  T_2208;
  wire  T_2211;
  reg [2:0] T_2219;
  reg [31:0] GEN_98;
  wire  T_2228;
  wire  T_2231;
  wire  T_2232;
  wire  T_2233;
  wire [2:0] T_2240_0;
  wire [2:0] T_2240_1;
  wire [2:0] T_2240_2;
  wire  T_2242;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  reg [2:0] T_2252;
  reg [31:0] GEN_99;
  wire  T_2254;
  wire [3:0] T_2256;
  wire [2:0] T_2257;
  wire [2:0] GEN_46;
  wire  T_2258;
  wire [2:0] T_2259;
  wire  T_2260;
  reg  T_2262;
  reg [31:0] GEN_100;
  wire  T_2264;
  wire  T_2265;
  wire [1:0] T_2267;
  wire  T_2268;
  wire  GEN_47;
  wire  T_2270;
  wire  T_2271;
  wire [1:0] T_2273;
  wire  T_2274;
  wire  GEN_48;
  wire  T_2276;
  wire  T_2280;
  wire  T_2282;
  wire  T_2283;
  wire [3:0] GEN_49;
  wire  T_2287;
  wire  T_2288;
  wire  T_2293;
  wire [2:0] T_2300_0;
  wire [2:0] T_2300_1;
  wire [2:0] T_2300_2;
  wire  T_2302;
  wire  T_2303;
  wire  T_2304;
  wire  T_2307;
  wire  T_2308;
  wire  T_2310;
  reg [2:0] T_2312;
  reg [31:0] GEN_101;
  wire  T_2314;
  wire [3:0] T_2316;
  wire [2:0] T_2317;
  wire [2:0] GEN_50;
  wire  T_2318;
  wire [2:0] T_2319;
  wire  T_2320;
  wire  T_2321;
  wire [3:0] GEN_452;
  wire  T_2324;
  wire  T_2325;
  wire  T_2326;
  wire  T_2327;
  wire [2:0] T_2335_0;
  wire [3:0] GEN_453;
  wire  T_2337;
  wire [1:0] T_2345_0;
  wire [1:0] T_2345_1;
  wire [3:0] GEN_454;
  wire  T_2347;
  wire [3:0] GEN_455;
  wire  T_2348;
  wire  T_2351;
  wire  T_2352;
  wire  T_2354;
  reg [2:0] T_2356;
  reg [31:0] GEN_102;
  wire  T_2358;
  wire [3:0] T_2360;
  wire [2:0] T_2361;
  wire [2:0] GEN_51;
  wire  T_2362;
  wire [2:0] T_2363;
  wire  T_2364;
  reg  T_2366;
  reg [31:0] GEN_103;
  wire  T_2368;
  wire  T_2369;
  wire [1:0] T_2371;
  wire  T_2372;
  wire  GEN_52;
  wire  T_2374;
  wire  T_2375;
  wire [1:0] T_2377;
  wire  T_2378;
  wire  GEN_53;
  wire  T_2380;
  wire  T_2382;
  wire  T_2383;
  wire [25:0] GEN_54;
  wire [3:0] GEN_55;
  wire  T_2386;
  wire [3:0] T_2392_0;
  wire [3:0] T_2392_1;
  wire  T_2394;
  wire  T_2395;
  wire  T_2398;
  wire  T_2400;
  wire  T_2401;
  wire  T_2403;
  wire  T_2404;
  wire  T_2405;
  wire  T_2407;
  wire  T_2408;
  wire  T_2411;
  wire  T_2412;
  wire  T_2414;
  wire  T_2415;
  wire [2:0] T_2422_0;
  wire [2:0] T_2422_1;
  wire [2:0] T_2422_2;
  wire  T_2424;
  wire  T_2425;
  wire  T_2426;
  wire  T_2429;
  wire  T_2430;
  wire  T_2433;
  wire  T_2435;
  wire  T_2436;
  wire  T_2437;
  wire  T_2438;
  wire [2:0] T_2445_0;
  wire [2:0] T_2445_1;
  wire [2:0] T_2445_2;
  wire  T_2447;
  wire  T_2448;
  wire  T_2449;
  wire  T_2452;
  wire  T_2453;
  wire [2:0] T_2461_0;
  wire [2:0] T_2461_1;
  wire [2:0] T_2461_2;
  wire  T_2463;
  wire  T_2464;
  wire  T_2465;
  wire  T_2468;
  wire  T_2469;
  wire  T_2470;
  wire [7:0] GEN_458;
  wire [8:0] T_2472;
  wire [7:0] T_2473;
  wire [7:0] T_2474;
  wire [7:0] T_2476;
  wire [7:0] T_2477;
  wire [7:0] T_2478;
  wire [7:0] T_2480;
  wire [2:0] GEN_56;
  wire  GEN_57;
  wire [1:0] GEN_58;
  wire [7:0] GEN_65;
  wire  T_2484;
  wire  T_2486;
  wire  T_2488;
  wire  T_2489;
  wire [2:0] T_2496_0;
  wire [2:0] T_2496_1;
  wire [2:0] T_2496_2;
  wire  T_2498;
  wire  T_2499;
  wire  T_2500;
  wire  T_2503;
  wire  T_2504;
  wire  T_2505;
  wire [7:0] GEN_460;
  wire [8:0] T_2507;
  wire [7:0] T_2508;
  wire [7:0] T_2509;
  wire [7:0] T_2513;
  wire [7:0] T_2514;
  wire [7:0] GEN_69;
  wire [2:0] GEN_75;
  wire  GEN_76;
  wire [1:0] GEN_77;
  wire [7:0] GEN_84;
  wire [3:0] T_2520_0;
  wire [3:0] T_2520_1;
  wire [3:0] T_2520_2;
  wire [3:0] T_2520_3;
  wire  T_2522;
  wire  T_2523;
  wire  T_2524;
  wire  T_2525;
  wire  T_2528;
  wire  T_2529;
  wire  T_2530;
  wire  T_2531;
  wire  T_2533;
  wire  T_2534;
  wire  T_2536;
  wire  T_2537;
  wire [2:0] T_2572_addr_beat;
  wire [25:0] T_2572_addr_block;
  wire [1:0] T_2572_client_xact_id;
  wire  T_2572_voluntary;
  wire [2:0] T_2572_r_type;
  wire [63:0] T_2572_data;
  wire  T_2572_client_id;
  wire [2:0] T_2639_addr_beat;
  wire [1:0] T_2639_client_xact_id;
  wire [2:0] T_2639_manager_xact_id;
  wire  T_2639_is_builtin_type;
  wire [3:0] T_2639_g_type;
  wire [63:0] T_2639_data;
  wire  T_2639_client_id;
  wire [3:0] T_2679_0;
  wire [3:0] T_2679_1;
  wire  T_2681;
  wire  T_2682;
  wire  T_2685;
  wire  T_2687;
  wire  T_2688;
  wire  T_2691;
  wire  T_2695;
  wire  T_2699;
  wire  T_2702;
  wire  T_2709;
  wire [2:0] T_2716_0;
  wire [2:0] T_2716_1;
  wire [2:0] T_2716_2;
  wire  T_2718;
  wire  T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [7:0] GEN_0;
  wire [7:0] GEN_88;
  wire [2:0] GEN_465;
  wire [7:0] GEN_89;
  wire [2:0] GEN_466;
  wire [7:0] GEN_90;
  wire [7:0] GEN_91;
  wire [7:0] GEN_92;
  wire [7:0] GEN_93;
  wire [7:0] GEN_94;
  wire  T_2726;
  wire [7:0] GEN_1;
  wire  T_2727;
  wire [7:0] GEN_2;
  wire  T_2728;
  wire [7:0] GEN_3;
  wire  T_2729;
  wire [7:0] GEN_4;
  wire  T_2730;
  wire [7:0] GEN_5;
  wire  T_2731;
  wire [7:0] GEN_6;
  wire  T_2732;
  wire [7:0] GEN_7;
  wire  T_2733;
  wire [7:0] GEN_488;
  wire [8:0] T_2735;
  wire [7:0] T_2736;
  wire [7:0] GEN_489;
  wire [8:0] T_2738;
  wire [7:0] T_2739;
  wire [7:0] GEN_490;
  wire [8:0] T_2741;
  wire [7:0] T_2742;
  wire [7:0] GEN_491;
  wire [8:0] T_2744;
  wire [7:0] T_2745;
  wire [7:0] GEN_492;
  wire [8:0] T_2747;
  wire [7:0] T_2748;
  wire [7:0] GEN_493;
  wire [8:0] T_2750;
  wire [7:0] T_2751;
  wire [7:0] GEN_494;
  wire [8:0] T_2753;
  wire [7:0] T_2754;
  wire [7:0] GEN_495;
  wire [8:0] T_2756;
  wire [7:0] T_2757;
  wire [7:0] T_2763_0;
  wire [7:0] T_2763_1;
  wire [7:0] T_2763_2;
  wire [7:0] T_2763_3;
  wire [7:0] T_2763_4;
  wire [7:0] T_2763_5;
  wire [7:0] T_2763_6;
  wire [7:0] T_2763_7;
  wire [15:0] T_2765;
  wire [15:0] T_2766;
  wire [31:0] T_2767;
  wire [15:0] T_2768;
  wire [15:0] T_2769;
  wire [31:0] T_2770;
  wire [63:0] T_2771;
  wire [63:0] T_2772;
  wire [63:0] T_2773;
  wire [63:0] GEN_8;
  wire [63:0] GEN_144;
  wire [63:0] GEN_145;
  wire [63:0] GEN_146;
  wire [63:0] GEN_147;
  wire [63:0] GEN_148;
  wire [63:0] GEN_149;
  wire [63:0] GEN_150;
  wire [63:0] T_2774;
  wire [63:0] T_2775;
  wire [63:0] GEN_9;
  wire [63:0] GEN_151;
  wire [63:0] GEN_152;
  wire [63:0] GEN_153;
  wire [63:0] GEN_154;
  wire [63:0] GEN_155;
  wire [63:0] GEN_156;
  wire [63:0] GEN_157;
  wire [63:0] GEN_158;
  wire [63:0] GEN_177;
  wire [63:0] GEN_178;
  wire [63:0] GEN_179;
  wire [63:0] GEN_180;
  wire [63:0] GEN_181;
  wire [63:0] GEN_182;
  wire [63:0] GEN_183;
  wire [63:0] GEN_184;
  wire [1:0] T_2806_state;
  wire  T_2832;
  wire  T_2833;
  wire [2:0] T_2839_0;
  wire [2:0] T_2839_1;
  wire [2:0] T_2839_2;
  wire  T_2841;
  wire  T_2842;
  wire  T_2843;
  wire  T_2846;
  wire  T_2847;
  wire  T_2848;
  wire [7:0] GEN_503;
  wire [8:0] T_2850;
  wire [7:0] T_2851;
  wire [7:0] T_2852;
  wire [7:0] T_2854;
  wire [7:0] T_2855;
  wire [7:0] T_2856;
  wire [7:0] T_2857;
  wire [2:0] T_2865_0;
  wire [2:0] T_2865_1;
  wire [2:0] T_2865_2;
  wire  T_2867;
  wire  T_2868;
  wire  T_2869;
  wire  T_2872;
  wire  T_2873;
  wire  T_2874;
  wire [7:0] GEN_505;
  wire [8:0] T_2877;
  wire [7:0] T_2878;
  wire [7:0] T_2881;
  wire [7:0] T_2882;
  wire [7:0] T_2883;
  wire [7:0] GEN_191;
  wire  GEN_193;
  wire  T_2893;
  wire [2:0] T_2900_0;
  wire [2:0] T_2900_1;
  wire [2:0] T_2900_2;
  wire  T_2902;
  wire  T_2903;
  wire  T_2904;
  wire  T_2907;
  wire  T_2908;
  wire  T_2910;
  reg [2:0] T_2912;
  reg [31:0] GEN_104;
  wire  T_2914;
  wire [3:0] T_2916;
  wire [2:0] T_2917;
  wire [2:0] GEN_194;
  wire  T_2918;
  wire [2:0] T_2919;
  wire  T_2920;
  wire  T_2923;
  wire  T_2924;
  wire  T_2925;
  wire [2:0] T_2933_0;
  wire [3:0] GEN_510;
  wire  T_2935;
  wire  T_2943_0;
  wire [3:0] GEN_511;
  wire  T_2945;
  wire  T_2948;
  wire  T_2950;
  reg [2:0] T_2952;
  reg [31:0] GEN_105;
  wire  T_2954;
  wire [3:0] T_2956;
  wire [2:0] T_2957;
  wire [2:0] GEN_195;
  wire  T_2958;
  wire [2:0] T_2959;
  wire  T_2960;
  reg  T_2962;
  reg [31:0] GEN_106;
  wire  T_2964;
  wire  T_2965;
  wire [1:0] T_2967;
  wire  T_2968;
  wire  GEN_196;
  wire  T_2970;
  wire  T_2971;
  wire [1:0] T_2973;
  wire  T_2974;
  wire  GEN_197;
  wire  T_2976;
  wire  T_2977;
  wire [2:0] T_2983_0;
  wire [2:0] T_2983_1;
  wire [2:0] T_2983_2;
  wire  T_2985;
  wire  T_2986;
  wire  T_2987;
  wire  T_2990;
  wire  T_2991;
  wire [7:0] T_2992;
  wire  T_2993;
  wire  T_2995;
  wire  T_2996;
  wire [1:0] T_3004_0;
  wire  T_3006;
  wire [2:0] T_3009;
  wire [2:0] T_3045_addr_beat;
  wire [25:0] T_3045_addr_block;
  wire [2:0] T_3045_client_xact_id;
  wire  T_3045_voluntary;
  wire [2:0] T_3045_r_type;
  wire [63:0] T_3045_data;
  wire [63:0] GEN_10;
  wire [63:0] GEN_198;
  wire [63:0] GEN_199;
  wire [63:0] GEN_200;
  wire [63:0] GEN_201;
  wire [63:0] GEN_202;
  wire [63:0] GEN_203;
  wire [63:0] GEN_204;
  wire  T_3074;
  wire  T_3076;
  wire [2:0] T_3087_0;
  wire  T_3089;
  wire  T_3092;
  wire  T_3093;
  reg [2:0] T_3095;
  reg [31:0] GEN_107;
  wire  T_3097;
  wire [3:0] T_3099;
  wire [2:0] T_3100;
  wire [2:0] GEN_205;
  wire  T_3101;
  wire [2:0] T_3102;
  wire  T_3103;
  wire  T_3109;
  wire  T_3110;
  wire [2:0] T_3118_0;
  wire [3:0] GEN_518;
  wire  T_3120;
  wire  T_3128_0;
  wire [3:0] GEN_519;
  wire  T_3130;
  wire  T_3133;
  wire  T_3135;
  reg [2:0] T_3137;
  reg [31:0] GEN_108;
  wire  T_3139;
  wire [3:0] T_3141;
  wire [2:0] T_3142;
  wire [2:0] GEN_206;
  wire  T_3143;
  wire [2:0] T_3144;
  wire  T_3145;
  reg  T_3147;
  reg [31:0] GEN_109;
  wire  T_3149;
  wire  T_3150;
  wire [1:0] T_3152;
  wire  T_3153;
  wire  GEN_207;
  wire  T_3155;
  wire  T_3156;
  wire [1:0] T_3158;
  wire  T_3159;
  wire  GEN_208;
  wire  T_3161;
  wire  T_3162;
  wire [7:0] T_3163;
  wire  T_3164;
  wire  T_3166;
  wire  T_3168;
  wire  T_3169;
  wire  T_3172;
  wire  T_3173;
  wire  T_3174;
  wire  T_3175;
  wire  T_3176;
  wire  T_3177;
  wire  T_3178;
  wire  T_3179;
  wire  T_3180;
  wire  T_3181;
  wire  T_3182;
  wire [5:0] T_3185;
  wire [25:0] T_3216_addr_block;
  wire [2:0] T_3216_client_xact_id;
  wire [2:0] T_3216_addr_beat;
  wire  T_3216_is_builtin_type;
  wire [2:0] T_3216_a_type;
  wire [11:0] T_3216_union;
  wire [63:0] T_3216_data;
  wire [7:0] GEN_11;
  wire [7:0] GEN_209;
  wire [7:0] GEN_210;
  wire [7:0] GEN_211;
  wire [7:0] GEN_212;
  wire [7:0] GEN_213;
  wire [7:0] GEN_214;
  wire [7:0] GEN_215;
  wire [5:0] T_3281;
  wire [5:0] T_3282;
  wire [11:0] T_3283;
  wire [7:0] T_3285;
  wire [8:0] T_3286;
  wire [8:0] T_3288;
  wire [5:0] T_3300;
  wire [5:0] T_3302;
  wire [11:0] T_3304;
  wire [11:0] T_3306;
  wire [11:0] T_3308;
  wire [11:0] T_3310;
  wire [11:0] T_3312;
  wire [25:0] T_3341_addr_block;
  wire [2:0] T_3341_client_xact_id;
  wire [2:0] T_3341_addr_beat;
  wire  T_3341_is_builtin_type;
  wire [2:0] T_3341_a_type;
  wire [11:0] T_3341_union;
  wire [63:0] T_3341_data;
  wire [63:0] GEN_12;
  wire [63:0] GEN_216;
  wire [63:0] GEN_217;
  wire [63:0] GEN_218;
  wire [63:0] GEN_219;
  wire [63:0] GEN_220;
  wire [63:0] GEN_221;
  wire [63:0] GEN_222;
  wire [25:0] T_3369_addr_block;
  wire [2:0] T_3369_client_xact_id;
  wire [2:0] T_3369_addr_beat;
  wire  T_3369_is_builtin_type;
  wire [2:0] T_3369_a_type;
  wire [11:0] T_3369_union;
  wire [63:0] T_3369_data;
  wire  T_3398;
  wire [3:0] GEN_223;
  wire [2:0] T_3408_0;
  wire [2:0] T_3408_1;
  wire [3:0] GEN_527;
  wire  T_3410;
  wire [3:0] GEN_528;
  wire  T_3411;
  wire  T_3414;
  wire  T_3420_0;
  wire [3:0] GEN_529;
  wire  T_3422;
  wire  T_3425;
  wire  T_3426;
  wire [7:0] GEN_13;
  wire [7:0] GEN_224;
  wire [7:0] GEN_225;
  wire [7:0] GEN_226;
  wire [7:0] GEN_227;
  wire [7:0] GEN_228;
  wire [7:0] GEN_229;
  wire [7:0] GEN_230;
  wire  T_3427;
  wire [7:0] GEN_14;
  wire  T_3428;
  wire [7:0] GEN_15;
  wire  T_3429;
  wire [7:0] GEN_16;
  wire  T_3430;
  wire [7:0] GEN_17;
  wire  T_3431;
  wire [7:0] GEN_18;
  wire  T_3432;
  wire [7:0] GEN_19;
  wire  T_3433;
  wire [7:0] GEN_20;
  wire  T_3434;
  wire [7:0] GEN_554;
  wire [8:0] T_3436;
  wire [7:0] T_3437;
  wire [7:0] GEN_555;
  wire [8:0] T_3439;
  wire [7:0] T_3440;
  wire [7:0] GEN_556;
  wire [8:0] T_3442;
  wire [7:0] T_3443;
  wire [7:0] GEN_557;
  wire [8:0] T_3445;
  wire [7:0] T_3446;
  wire [7:0] GEN_558;
  wire [8:0] T_3448;
  wire [7:0] T_3449;
  wire [7:0] GEN_559;
  wire [8:0] T_3451;
  wire [7:0] T_3452;
  wire [7:0] GEN_560;
  wire [8:0] T_3454;
  wire [7:0] T_3455;
  wire [7:0] GEN_561;
  wire [8:0] T_3457;
  wire [7:0] T_3458;
  wire [7:0] T_3464_0;
  wire [7:0] T_3464_1;
  wire [7:0] T_3464_2;
  wire [7:0] T_3464_3;
  wire [7:0] T_3464_4;
  wire [7:0] T_3464_5;
  wire [7:0] T_3464_6;
  wire [7:0] T_3464_7;
  wire [15:0] T_3466;
  wire [15:0] T_3467;
  wire [31:0] T_3468;
  wire [15:0] T_3469;
  wire [15:0] T_3470;
  wire [31:0] T_3471;
  wire [63:0] T_3472;
  wire [63:0] T_3473;
  wire [63:0] T_3474;
  wire [63:0] GEN_21;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [63:0] GEN_286;
  wire [63:0] T_3475;
  wire [63:0] T_3476;
  wire [63:0] GEN_22;
  wire [63:0] GEN_287;
  wire [63:0] GEN_288;
  wire [63:0] GEN_289;
  wire [63:0] GEN_290;
  wire [63:0] GEN_291;
  wire [63:0] GEN_292;
  wire [63:0] GEN_293;
  wire [63:0] GEN_294;
  wire [63:0] GEN_313;
  wire [63:0] GEN_314;
  wire [63:0] GEN_315;
  wire [63:0] GEN_316;
  wire [63:0] GEN_317;
  wire [63:0] GEN_318;
  wire [63:0] GEN_319;
  wire [63:0] GEN_320;
  wire  T_3477;
  wire  T_3478;
  wire  T_3489;
  wire  T_3491;
  wire [2:0] T_3499_0;
  wire [3:0] GEN_570;
  wire  T_3501;
  wire [1:0] T_3509_0;
  wire [1:0] T_3509_1;
  wire [3:0] GEN_571;
  wire  T_3511;
  wire [3:0] GEN_572;
  wire  T_3512;
  wire  T_3515;
  wire  T_3516;
  wire  T_3518;
  reg [2:0] T_3520;
  reg [31:0] GEN_110;
  wire  T_3522;
  wire [3:0] T_3524;
  wire [2:0] T_3525;
  wire [2:0] GEN_321;
  wire  T_3526;
  wire [2:0] T_3527;
  wire  T_3528;
  wire  T_3529;
  reg [2:0] T_3535;
  reg [31:0] GEN_111;
  reg  T_3545;
  reg [31:0] GEN_112;
  wire  T_3547;
  wire  T_3548;
  wire [1:0] T_3550;
  wire  T_3551;
  wire  GEN_323;
  wire  T_3553;
  wire  T_3554;
  wire [1:0] T_3556;
  wire  T_3557;
  wire  GEN_324;
  wire  T_3559;
  wire  T_3564;
  wire [2:0] T_3573_0;
  wire [2:0] T_3573_1;
  wire [3:0] GEN_575;
  wire  T_3575;
  wire [3:0] GEN_576;
  wire  T_3576;
  wire  T_3579;
  wire [1:0] T_3585_0;
  wire [1:0] T_3585_1;
  wire [3:0] GEN_577;
  wire  T_3587;
  wire [3:0] GEN_578;
  wire  T_3588;
  wire  T_3591;
  wire  T_3592;
  wire  T_3593;
  wire [7:0] GEN_579;
  wire [8:0] T_3595;
  wire [7:0] T_3596;
  wire [7:0] T_3597;
  wire [7:0] T_3599;
  wire [7:0] T_3600;
  wire [7:0] T_3601;
  wire [7:0] T_3602;
  wire [2:0] T_3610_0;
  wire [2:0] T_3610_1;
  wire [2:0] T_3610_2;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3617;
  wire  T_3618;
  wire  T_3619;
  wire [7:0] GEN_581;
  wire [8:0] T_3622;
  wire [7:0] T_3623;
  wire [7:0] T_3626;
  wire [7:0] T_3627;
  wire [2:0] T_3637_0;
  wire [2:0] T_3637_1;
  wire [3:0] GEN_583;
  wire  T_3639;
  wire [3:0] GEN_584;
  wire  T_3640;
  wire  T_3643;
  wire  T_3649_0;
  wire [3:0] GEN_585;
  wire  T_3651;
  wire  T_3654;
  wire  T_3655;
  wire [7:0] GEN_586;
  wire [8:0] T_3658;
  wire [7:0] T_3659;
  wire [7:0] T_3661;
  wire [7:0] T_3662;
  wire [7:0] T_3663;
  wire [7:0] T_3664;
  wire [7:0] GEN_335;
  wire  T_3666;
  wire  T_3667;
  wire  T_3670;
  wire  T_3672;
  wire  T_3689;
  wire [2:0] T_3690;
  wire  T_3691;
  wire [2:0] T_3692;
  wire  T_3693;
  wire [2:0] T_3694;
  wire  T_3695;
  wire [2:0] T_3696;
  wire  T_3697;
  wire [2:0] T_3698;
  wire  T_3699;
  wire [2:0] T_3700;
  wire  T_3701;
  wire [2:0] T_3702;
  wire  T_3703;
  wire [1:0] T_3708;
  wire [2:0] T_3709;
  wire [2:0] T_3741_addr_beat;
  wire [1:0] T_3741_client_xact_id;
  wire [2:0] T_3741_manager_xact_id;
  wire  T_3741_is_builtin_type;
  wire [3:0] T_3741_g_type;
  wire [63:0] T_3741_data;
  wire  T_3741_client_id;
  wire [63:0] GEN_23;
  wire [63:0] GEN_336;
  wire [63:0] GEN_337;
  wire [63:0] GEN_338;
  wire [63:0] GEN_339;
  wire [63:0] GEN_340;
  wire [63:0] GEN_341;
  wire [63:0] GEN_342;
  wire [2:0] T_3780_0;
  wire [3:0] GEN_594;
  wire  T_3782;
  wire [1:0] T_3790_0;
  wire [1:0] T_3790_1;
  wire [3:0] GEN_595;
  wire  T_3792;
  wire [3:0] GEN_596;
  wire  T_3793;
  wire  T_3796;
  wire  T_3797;
  wire  T_3799;
  reg [2:0] T_3801;
  reg [31:0] GEN_113;
  wire  T_3803;
  wire [3:0] T_3805;
  wire [2:0] T_3806;
  wire [2:0] GEN_343;
  wire  T_3807;
  wire [2:0] T_3808;
  wire  T_3809;
  wire  T_3814;
  wire  T_3816;
  wire [2:0] T_3824_0;
  wire [2:0] T_3824_1;
  wire [3:0] GEN_598;
  wire  T_3826;
  wire [3:0] GEN_599;
  wire  T_3827;
  wire  T_3830;
  wire [1:0] T_3836_0;
  wire [1:0] T_3836_1;
  wire [3:0] GEN_600;
  wire  T_3838;
  wire [3:0] GEN_601;
  wire  T_3839;
  wire  T_3842;
  wire  T_3843;
  wire [7:0] T_3844;
  wire  T_3845;
  wire  T_3846;
  wire  T_3847;
  wire  GEN_348;
  wire  GEN_349;
  wire [2:0] GEN_350;
  wire [1:0] GEN_351;
  wire [2:0] GEN_352;
  wire  GEN_353;
  wire [3:0] GEN_354;
  wire [63:0] GEN_355;
  wire  GEN_356;
  wire  GEN_361;
  wire  T_3854;
  wire [1:0] GEN_362;
  wire [2:0] T_3869_0;
  wire  T_3871;
  wire  T_3874;
  wire  T_3875;
  wire  T_3876;
  wire  T_3879;
  wire  T_3881;
  wire  T_3882;
  wire [2:0] T_3892_0;
  wire [2:0] T_3892_1;
  wire [2:0] T_3892_2;
  wire  T_3894;
  wire  T_3895;
  wire  T_3896;
  wire  T_3899;
  wire  T_3900;
  wire  T_3901;
  wire  T_3902;
  wire  T_3903;
  wire  T_3905;
  wire  T_3906;
  wire [8:0] T_3910;
  wire [7:0] T_3911;
  wire [7:0] T_3917_0;
  wire  T_3925;
  wire [7:0] T_3926;
  wire [7:0] T_3928;
  wire [7:0] T_3929;
  wire  T_3930;
  wire  T_3931;
  wire  T_3932;
  wire  T_3933;
  wire  T_3934;
  wire  T_3935;
  wire  T_3936;
  wire  T_3937;
  wire [7:0] GEN_603;
  wire [8:0] T_3939;
  wire [7:0] T_3940;
  wire [7:0] GEN_604;
  wire [8:0] T_3942;
  wire [7:0] T_3943;
  wire [7:0] GEN_605;
  wire [8:0] T_3945;
  wire [7:0] T_3946;
  wire [7:0] GEN_606;
  wire [8:0] T_3948;
  wire [7:0] T_3949;
  wire [7:0] GEN_607;
  wire [8:0] T_3951;
  wire [7:0] T_3952;
  wire [7:0] GEN_608;
  wire [8:0] T_3954;
  wire [7:0] T_3955;
  wire [7:0] GEN_609;
  wire [8:0] T_3957;
  wire [7:0] T_3958;
  wire [7:0] GEN_610;
  wire [8:0] T_3960;
  wire [7:0] T_3961;
  wire [7:0] T_3967_0;
  wire [7:0] T_3967_1;
  wire [7:0] T_3967_2;
  wire [7:0] T_3967_3;
  wire [7:0] T_3967_4;
  wire [7:0] T_3967_5;
  wire [7:0] T_3967_6;
  wire [7:0] T_3967_7;
  wire [15:0] T_3969;
  wire [15:0] T_3970;
  wire [31:0] T_3971;
  wire [15:0] T_3972;
  wire [15:0] T_3973;
  wire [31:0] T_3974;
  wire [63:0] T_3975;
  wire [63:0] T_3976;
  wire [63:0] GEN_24;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [63:0] GEN_366;
  wire [63:0] GEN_367;
  wire [63:0] GEN_368;
  wire [63:0] GEN_369;
  wire [63:0] T_3977;
  wire [63:0] T_3978;
  wire [63:0] T_3979;
  wire [63:0] GEN_25;
  wire [63:0] GEN_370;
  wire [63:0] GEN_371;
  wire [63:0] GEN_372;
  wire [63:0] GEN_373;
  wire [63:0] GEN_374;
  wire [63:0] GEN_375;
  wire [63:0] GEN_376;
  wire [63:0] GEN_377;
  wire [7:0] T_3993_0;
  wire [7:0] T_4005;
  wire [7:0] GEN_26;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [7:0] GEN_381;
  wire [7:0] GEN_382;
  wire [7:0] GEN_383;
  wire [7:0] GEN_384;
  wire [7:0] T_4006;
  wire [7:0] GEN_27;
  wire [7:0] GEN_385;
  wire [7:0] GEN_386;
  wire [7:0] GEN_387;
  wire [7:0] GEN_388;
  wire [7:0] GEN_389;
  wire [7:0] GEN_390;
  wire [7:0] GEN_391;
  wire [7:0] GEN_392;
  wire [63:0] GEN_404;
  wire [63:0] GEN_405;
  wire [63:0] GEN_406;
  wire [63:0] GEN_407;
  wire [63:0] GEN_408;
  wire [63:0] GEN_409;
  wire [63:0] GEN_410;
  wire [63:0] GEN_411;
  wire [7:0] GEN_415;
  wire [7:0] GEN_416;
  wire [7:0] GEN_417;
  wire [7:0] GEN_418;
  wire [7:0] GEN_419;
  wire [7:0] GEN_420;
  wire [7:0] GEN_421;
  wire [7:0] GEN_422;
  wire  T_4009;
  wire  T_4010;
  wire  T_4011;
  wire  T_4012;
  wire  T_4013;
  wire  T_4014;
  wire  T_4015;
  wire  T_4017;
  wire  T_4019;
  wire [3:0] GEN_423;
  wire [7:0] GEN_424;
  wire [7:0] GEN_425;
  wire [7:0] GEN_426;
  wire [7:0] GEN_427;
  wire [7:0] GEN_428;
  wire [7:0] GEN_429;
  wire [7:0] GEN_430;
  wire [7:0] GEN_431;
  reg  GEN_28;
  reg [31:0] GEN_114;
  reg  GEN_29;
  reg [31:0] GEN_115;
  Queue_11 Queue_13_1 (
    .clk(Queue_13_1_clk),
    .reset(Queue_13_1_reset),
    .io_enq_ready(Queue_13_1_io_enq_ready),
    .io_enq_valid(Queue_13_1_io_enq_valid),
    .io_enq_bits_client_xact_id(Queue_13_1_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(Queue_13_1_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(Queue_13_1_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(Queue_13_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(Queue_13_1_io_enq_bits_a_type),
    .io_deq_ready(Queue_13_1_io_deq_ready),
    .io_deq_valid(Queue_13_1_io_deq_valid),
    .io_deq_bits_client_xact_id(Queue_13_1_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(Queue_13_1_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(Queue_13_1_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(Queue_13_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(Queue_13_1_io_deq_bits_a_type),
    .io_count(Queue_13_1_io_count)
  );
  assign io_inner_acquire_ready = T_2099;
  assign io_inner_grant_valid = GEN_361;
  assign io_inner_grant_bits_addr_beat = GEN_350;
  assign io_inner_grant_bits_client_xact_id = GEN_351;
  assign io_inner_grant_bits_manager_xact_id = GEN_352;
  assign io_inner_grant_bits_is_builtin_type = GEN_353;
  assign io_inner_grant_bits_g_type = GEN_354;
  assign io_inner_grant_bits_data = GEN_355;
  assign io_inner_grant_bits_client_id = GEN_356;
  assign io_inner_finish_ready = T_2977;
  assign io_inner_probe_valid = T_2211;
  assign io_inner_probe_bits_addr_block = T_2155_addr_block;
  assign io_inner_probe_bits_p_type = T_2155_p_type;
  assign io_inner_probe_bits_client_id = T_2155_client_id;
  assign io_inner_release_ready = T_2709;
  assign io_outer_acquire_valid = T_3169;
  assign io_outer_acquire_bits_addr_block = T_3369_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3369_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3369_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3369_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3369_a_type;
  assign io_outer_acquire_bits_union = T_3369_union;
  assign io_outer_acquire_bits_data = T_3369_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2996;
  assign io_outer_release_bits_addr_beat = T_3045_addr_beat;
  assign io_outer_release_bits_addr_block = T_3045_addr_block;
  assign io_outer_release_bits_client_xact_id = T_3045_client_xact_id;
  assign io_outer_release_bits_voluntary = T_3045_voluntary;
  assign io_outer_release_bits_r_type = T_3045_r_type;
  assign io_outer_release_bits_data = T_3045_data;
  assign io_outer_grant_ready = T_2977;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_28;
  assign io_outer_finish_bits_manager_id = GEN_29;
  assign io_alloc_iacq_matches = T_1842;
  assign io_alloc_iacq_can = T_1733;
  assign io_alloc_irel_matches = T_1845;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1848;
  assign io_alloc_oprb_can = 1'h0;
  assign T_44 = T_4017;
  assign T_69 = T_99_addr_beat;
  assign T_99_client_xact_id = T_1930_client_xact_id;
  assign T_99_addr_beat = T_1930_addr_beat;
  assign T_99_client_id = T_1930_client_id;
  assign T_99_is_builtin_type = T_1930_is_builtin_type;
  assign T_99_a_type = T_1930_a_type;
  assign T_144_pending = T_2380;
  assign T_144_up_idx = T_2319;
  assign T_144_up_done = T_2320;
  assign T_144_down_idx = T_2363;
  assign T_144_down_done = T_2364;
  assign T_153 = T_1960;
  assign T_155 = T_3808;
  assign T_157 = T_3809;
  assign T_166_pending = T_3559;
  assign T_166_up_idx = T_3527;
  assign T_166_up_done = T_3528;
  assign T_166_down_idx = 3'h0;
  assign T_166_down_done = T_3529;
  assign T_186_pending = T_3161;
  assign T_186_up_idx = T_3102;
  assign T_186_up_done = T_3103;
  assign T_186_down_idx = T_3144;
  assign T_186_down_done = T_3145;
  assign T_210_pending = T_2976;
  assign T_210_up_idx = T_2919;
  assign T_210_up_done = T_2920;
  assign T_210_down_idx = T_2959;
  assign T_210_down_done = T_2960;
  assign GEN_432 = {{7'd0}, 1'h0};
  assign T_219 = T_201 != GEN_432;
  assign T_220 = T_199 | T_219;
  assign T_221 = T_220 | T_210_pending;
  assign T_247_sharers = 1'h0;
  assign T_299_state = {{1'd0}, 1'h0};
  assign T_395_inner_sharers = T_247_sharers;
  assign T_395_outer_state = T_299_state;
  assign T_1733 = T_55 == 4'h0;
  assign T_1734 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1735 = T_1733 & T_1734;
  assign T_1736 = T_1735 & io_alloc_iacq_should;
  assign T_1745_0 = 3'h3;
  assign T_1747 = T_1745_0 == io_inner_acquire_bits_a_type;
  assign T_1750 = io_inner_acquire_bits_is_builtin_type & T_1747;
  assign T_1751 = T_1736 & T_1750;
  assign T_1760_0 = 3'h3;
  assign T_1762 = T_1760_0 == io_inner_acquire_bits_a_type;
  assign T_1765 = io_inner_acquire_bits_is_builtin_type & T_1762;
  assign T_1767 = T_1765 == 1'h0;
  assign GEN_433 = {{2'd0}, 1'h0};
  assign T_1769 = io_inner_acquire_bits_addr_beat == GEN_433;
  assign T_1770 = T_1767 | T_1769;
  assign T_1772 = T_1770 == 1'h0;
  assign T_1773 = T_1751 & T_1772;
  assign T_1775 = T_1773 == 1'h0;
  assign T_1776 = T_1775 | reset;
  assign T_1778 = T_1776 == 1'h0;
  assign T_1779 = T_55 != 4'h0;
  assign T_1780 = T_1779 & T_153;
  assign T_1782 = T_99_a_type == 3'h5;
  assign T_1784 = T_99_a_type == 3'h6;
  assign T_1785 = T_1782 | T_1784;
  assign T_1786 = T_99_is_builtin_type & T_1785;
  assign T_1787 = T_1780 & T_1786;
  assign T_1789 = T_1787 == 1'h0;
  assign T_1790 = T_1789 | reset;
  assign T_1792 = T_1790 == 1'h0;
  assign T_1796 = T_99_a_type == 3'h4;
  assign T_1797 = T_99_is_builtin_type & T_1796;
  assign T_1798 = T_1780 & T_1797;
  assign T_1800 = T_1798 == 1'h0;
  assign T_1801 = T_1800 | reset;
  assign T_1803 = T_1801 == 1'h0;
  assign T_1817_0 = 64'h0;
  assign T_1817_1 = 64'h0;
  assign T_1817_2 = 64'h0;
  assign T_1817_3 = 64'h0;
  assign T_1817_4 = 64'h0;
  assign T_1817_5 = 64'h0;
  assign T_1817_6 = 64'h0;
  assign T_1817_7 = 64'h0;
  assign T_1835_0 = 8'h0;
  assign T_1835_1 = 8'h0;
  assign T_1835_2 = 8'h0;
  assign T_1835_3 = 8'h0;
  assign T_1835_4 = 8'h0;
  assign T_1835_5 = 8'h0;
  assign T_1835_6 = 8'h0;
  assign T_1835_7 = 8'h0;
  assign T_1841 = io_inner_acquire_bits_addr_block == T_57;
  assign T_1842 = T_1779 & T_1841;
  assign T_1844 = io_inner_release_bits_addr_block == T_57;
  assign T_1845 = T_1779 & T_1844;
  assign T_1847 = io_outer_probe_bits_addr_block == T_57;
  assign T_1848 = T_1779 & T_1847;
  assign Queue_13_1_clk = clk;
  assign Queue_13_1_reset = reset;
  assign Queue_13_1_io_enq_valid = T_1929;
  assign Queue_13_1_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign Queue_13_1_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign Queue_13_1_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign Queue_13_1_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign Queue_13_1_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign Queue_13_1_io_deq_ready = GEN_349;
  assign T_1884 = T_1733 & io_alloc_iacq_should;
  assign T_1885 = T_1884 & io_inner_acquire_valid;
  assign T_1887 = T_99_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1896_0 = 3'h3;
  assign T_1898 = T_1896_0 == T_99_a_type;
  assign T_1901 = T_99_is_builtin_type & T_1898;
  assign T_1902 = T_1887 & T_1901;
  assign T_1903 = T_1902 & T_153;
  assign T_1904 = T_175 >> io_inner_acquire_bits_addr_beat;
  assign T_1905 = T_1904[0];
  assign T_1906 = T_1903 & T_1905;
  assign T_1908 = T_1906 & io_inner_acquire_valid;
  assign T_1917_0 = 3'h3;
  assign T_1919 = T_1917_0 == io_inner_acquire_bits_a_type;
  assign T_1922 = io_inner_acquire_bits_is_builtin_type & T_1919;
  assign T_1924 = T_1922 == 1'h0;
  assign T_1927 = T_1924 | T_1769;
  assign T_1928 = T_1908 & T_1927;
  assign T_1929 = T_1885 | T_1928;
  assign T_1930_client_xact_id = Queue_13_1_io_deq_valid ? Queue_13_1_io_deq_bits_client_xact_id : Queue_13_1_io_enq_bits_client_xact_id;
  assign T_1930_addr_beat = Queue_13_1_io_deq_valid ? Queue_13_1_io_deq_bits_addr_beat : Queue_13_1_io_enq_bits_addr_beat;
  assign T_1930_client_id = Queue_13_1_io_deq_valid ? Queue_13_1_io_deq_bits_client_id : Queue_13_1_io_enq_bits_client_id;
  assign T_1930_is_builtin_type = Queue_13_1_io_deq_valid ? Queue_13_1_io_deq_bits_is_builtin_type : Queue_13_1_io_enq_bits_is_builtin_type;
  assign T_1930_a_type = Queue_13_1_io_deq_valid ? Queue_13_1_io_deq_bits_a_type : Queue_13_1_io_enq_bits_a_type;
  assign GEN_435 = {{1'd0}, 1'h0};
  assign T_1960 = Queue_13_1_io_count > GEN_435;
  assign T_1962 = T_1779 | io_alloc_iacq_should;
  assign T_1972_0 = 3'h2;
  assign T_1972_1 = 3'h3;
  assign T_1972_2 = 3'h4;
  assign T_1974 = T_1972_0 == io_inner_acquire_bits_a_type;
  assign T_1975 = T_1972_1 == io_inner_acquire_bits_a_type;
  assign T_1976 = T_1972_2 == io_inner_acquire_bits_a_type;
  assign T_1979 = T_1974 | T_1975;
  assign T_1980 = T_1979 | T_1976;
  assign T_1981 = io_inner_acquire_bits_is_builtin_type & T_1980;
  assign T_1982 = T_1734 & T_1981;
  assign GEN_436 = {{7'd0}, T_1982};
  assign T_1984 = 8'h0 - GEN_436;
  assign T_1985 = T_1984[7:0];
  assign T_1986 = ~ T_1985;
  assign GEN_437 = {{7'd0}, 1'h1};
  assign T_1988 = GEN_437 << io_inner_acquire_bits_addr_beat;
  assign T_1989 = ~ T_1988;
  assign T_1990 = T_1986 | T_1989;
  assign T_1991 = T_175 & T_1990;
  assign T_2001_0 = 3'h3;
  assign T_2003 = T_2001_0 == io_inner_acquire_bits_a_type;
  assign T_2006 = io_inner_acquire_bits_is_builtin_type & T_2003;
  assign T_2007 = T_1734 & T_2006;
  assign T_2010 = T_2007 & T_1769;
  assign T_2019 = T_2010 ? 8'hfe : 8'h0;
  assign T_2020 = T_1991 | T_2019;
  assign GEN_32 = T_1962 ? T_2020 : T_175;
  assign GEN_439 = {{3'd0}, 1'h0};
  assign T_2028 = 4'h8 * GEN_439;
  assign T_2030 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_2031 = io_inner_acquire_bits_is_builtin_type & T_2030;
  assign T_2033 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_2034 = io_inner_acquire_bits_is_builtin_type & T_2033;
  assign T_2035 = T_2031 | T_2034;
  assign T_2036 = io_inner_acquire_bits_union[5:1];
  assign T_2037 = T_2035 ? 5'h1 : T_2036;
  assign T_2038 = io_inner_acquire_bits_union[11:9];
  assign T_2039 = io_inner_acquire_bits_union[8:6];
  assign T_2052_0 = 3'h2;
  assign T_2052_1 = 3'h3;
  assign T_2052_2 = 3'h4;
  assign T_2054 = T_2052_0 == io_inner_acquire_bits_a_type;
  assign T_2055 = T_2052_1 == io_inner_acquire_bits_a_type;
  assign T_2056 = T_2052_2 == io_inner_acquire_bits_a_type;
  assign T_2059 = T_2054 | T_2055;
  assign T_2060 = T_2059 | T_2056;
  assign T_2061 = io_inner_acquire_bits_is_builtin_type & T_2060;
  assign T_2062 = T_1734 & T_2061;
  assign GEN_440 = {{7'd0}, T_2062};
  assign T_2064 = 8'h0 - GEN_440;
  assign T_2065 = T_2064[7:0];
  assign T_2066 = ~ T_2065;
  assign T_2070 = T_2066 | T_1989;
  assign T_2072 = T_2034 ? T_2070 : {{7'd0}, 1'h0};
  assign GEN_33 = T_1885 ? io_inner_acquire_bits_addr_block : T_57;
  assign GEN_34 = T_1885 ? 1'h0 : T_59;
  assign GEN_35 = T_1885 ? T_2028 : T_61;
  assign GEN_36 = T_1885 ? T_2037 : T_63;
  assign GEN_37 = T_1885 ? T_2038 : T_65;
  assign GEN_38 = T_1885 ? T_2039 : T_67;
  assign GEN_42 = T_1885 ? T_2072 : GEN_32;
  assign GEN_43 = T_1885 ? {{7'd0}, 1'h0} : T_177;
  assign GEN_44 = T_1885 ? 4'h5 : T_55;
  assign T_2075 = T_175 != GEN_432;
  assign T_2088_0 = 3'h3;
  assign T_2090 = T_2088_0 == T_99_a_type;
  assign T_2093 = T_99_is_builtin_type & T_2090;
  assign T_2094 = T_1887 & T_2093;
  assign T_2095 = T_2094 & T_153;
  assign T_2098 = T_2095 & T_1905;
  assign T_2099 = T_1733 | T_2098;
  assign T_2100 = ~ T_177;
  assign skip_outer_acquire = T_2100 == GEN_432;
  assign T_2109 = 3'h4 == T_99_a_type;
  assign T_2110 = T_2109 ? 2'h0 : 2'h2;
  assign T_2111 = 3'h6 == T_99_a_type;
  assign T_2112 = T_2111 ? 2'h0 : T_2110;
  assign T_2113 = 3'h5 == T_99_a_type;
  assign T_2114 = T_2113 ? 2'h2 : T_2112;
  assign T_2115 = 3'h2 == T_99_a_type;
  assign T_2116 = T_2115 ? 2'h0 : T_2114;
  assign T_2117 = 3'h0 == T_99_a_type;
  assign T_2118 = T_2117 ? 2'h2 : T_2116;
  assign T_2119 = 3'h3 == T_99_a_type;
  assign T_2120 = T_2119 ? 2'h0 : T_2118;
  assign T_2121 = 3'h1 == T_99_a_type;
  assign T_2122 = T_2121 ? 2'h2 : T_2120;
  assign GEN_444 = {{2'd0}, 1'h1};
  assign T_2123 = GEN_444 == T_99_a_type;
  assign T_2124 = T_2123 ? 2'h0 : 2'h2;
  assign T_2125 = GEN_433 == T_99_a_type;
  assign T_2126 = T_2125 ? 2'h1 : T_2124;
  assign T_2127 = T_99_is_builtin_type ? T_2122 : T_2126;
  assign T_2155_addr_block = T_57;
  assign T_2155_p_type = T_2127;
  assign T_2155_client_id = 1'h0;
  assign T_2183 = skip_outer_acquire == 1'h0;
  assign T_2184 = T_2183 ? 4'h6 : 4'h7;
  assign T_2193_pending = T_2276;
  assign T_2193_up_idx = 3'h0;
  assign T_2193_up_done = T_2201;
  assign T_2193_down_idx = T_2259;
  assign T_2193_down_done = T_2260;
  assign T_2201 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2202 = ~ T_2201;
  assign GEN_446 = {{1'd0}, 1'h1};
  assign T_2204 = GEN_446 << io_inner_probe_bits_client_id;
  assign T_2205 = ~ T_2204;
  assign GEN_447 = {{1'd0}, T_2202};
  assign T_2206 = GEN_447 | T_2205;
  assign GEN_448 = {{1'd0}, T_195};
  assign T_2207 = GEN_448 & T_2206;
  assign T_2208 = T_55 == 4'h5;
  assign T_2211 = T_2208 & T_195;
  assign T_2228 = io_inner_release_ready & io_inner_release_valid;
  assign T_2231 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2232 = T_1779 & T_2231;
  assign T_2233 = T_2228 & T_2232;
  assign T_2240_0 = 3'h0;
  assign T_2240_1 = 3'h1;
  assign T_2240_2 = 3'h2;
  assign T_2242 = T_2240_0 == io_inner_release_bits_r_type;
  assign T_2243 = T_2240_1 == io_inner_release_bits_r_type;
  assign T_2244 = T_2240_2 == io_inner_release_bits_r_type;
  assign T_2247 = T_2242 | T_2243;
  assign T_2248 = T_2247 | T_2244;
  assign T_2250 = T_2233 & T_2248;
  assign T_2254 = T_2252 == 3'h7;
  assign T_2256 = T_2252 + GEN_444;
  assign T_2257 = T_2256[2:0];
  assign GEN_46 = T_2250 ? T_2257 : T_2252;
  assign T_2258 = T_2250 & T_2254;
  assign T_2259 = T_2248 ? T_2252 : {{2'd0}, 1'h0};
  assign T_2260 = T_2248 ? T_2258 : T_2233;
  assign T_2264 = T_2260 == 1'h0;
  assign T_2265 = T_2201 & T_2264;
  assign T_2267 = T_2262 + 1'h1;
  assign T_2268 = T_2267[0:0];
  assign GEN_47 = T_2265 ? T_2268 : T_2262;
  assign T_2270 = T_2201 == 1'h0;
  assign T_2271 = T_2260 & T_2270;
  assign T_2273 = T_2262 - 1'h1;
  assign T_2274 = T_2273[0:0];
  assign GEN_48 = T_2271 ? T_2274 : GEN_47;
  assign T_2276 = T_2262 > 1'h0;
  assign T_2280 = T_195 | T_2193_pending;
  assign T_2282 = T_2280 == 1'h0;
  assign T_2283 = T_2208 & T_2282;
  assign GEN_49 = T_2283 ? T_2184 : GEN_44;
  assign T_2287 = T_1733 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2288 = T_2287 & io_inner_release_bits_voluntary;
  assign T_2293 = T_2228 & T_2288;
  assign T_2300_0 = 3'h0;
  assign T_2300_1 = 3'h1;
  assign T_2300_2 = 3'h2;
  assign T_2302 = T_2300_0 == io_inner_release_bits_r_type;
  assign T_2303 = T_2300_1 == io_inner_release_bits_r_type;
  assign T_2304 = T_2300_2 == io_inner_release_bits_r_type;
  assign T_2307 = T_2302 | T_2303;
  assign T_2308 = T_2307 | T_2304;
  assign T_2310 = T_2293 & T_2308;
  assign T_2314 = T_2312 == 3'h7;
  assign T_2316 = T_2312 + GEN_444;
  assign T_2317 = T_2316[2:0];
  assign GEN_50 = T_2310 ? T_2317 : T_2312;
  assign T_2318 = T_2310 & T_2314;
  assign T_2319 = T_2308 ? T_2312 : {{2'd0}, 1'h0};
  assign T_2320 = T_2308 ? T_2318 : T_2293;
  assign T_2321 = io_inner_grant_ready & io_inner_grant_valid;
  assign GEN_452 = {{1'd0}, 3'h0};
  assign T_2324 = io_inner_grant_bits_g_type == GEN_452;
  assign T_2325 = io_inner_grant_bits_is_builtin_type & T_2324;
  assign T_2326 = T_1779 & T_2325;
  assign T_2327 = T_2321 & T_2326;
  assign T_2335_0 = 3'h5;
  assign GEN_453 = {{1'd0}, T_2335_0};
  assign T_2337 = GEN_453 == io_inner_grant_bits_g_type;
  assign T_2345_0 = 2'h0;
  assign T_2345_1 = 2'h1;
  assign GEN_454 = {{2'd0}, T_2345_0};
  assign T_2347 = GEN_454 == io_inner_grant_bits_g_type;
  assign GEN_455 = {{2'd0}, T_2345_1};
  assign T_2348 = GEN_455 == io_inner_grant_bits_g_type;
  assign T_2351 = T_2347 | T_2348;
  assign T_2352 = io_inner_grant_bits_is_builtin_type ? T_2337 : T_2351;
  assign T_2354 = T_2327 & T_2352;
  assign T_2358 = T_2356 == 3'h7;
  assign T_2360 = T_2356 + GEN_444;
  assign T_2361 = T_2360[2:0];
  assign GEN_51 = T_2354 ? T_2361 : T_2356;
  assign T_2362 = T_2354 & T_2358;
  assign T_2363 = T_2352 ? T_2356 : {{2'd0}, 1'h0};
  assign T_2364 = T_2352 ? T_2362 : T_2327;
  assign T_2368 = T_2364 == 1'h0;
  assign T_2369 = T_2320 & T_2368;
  assign T_2371 = T_2366 + 1'h1;
  assign T_2372 = T_2371[0:0];
  assign GEN_52 = T_2369 ? T_2372 : T_2366;
  assign T_2374 = T_2320 == 1'h0;
  assign T_2375 = T_2364 & T_2374;
  assign T_2377 = T_2366 - 1'h1;
  assign T_2378 = T_2377[0:0];
  assign GEN_53 = T_2375 ? T_2378 : GEN_52;
  assign T_2380 = T_2366 > 1'h0;
  assign T_2382 = T_1733 & io_alloc_irel_should;
  assign T_2383 = T_2382 & io_inner_release_valid;
  assign GEN_54 = T_2383 ? io_inner_release_bits_addr_block : GEN_33;
  assign GEN_55 = T_2383 ? 4'h7 : GEN_49;
  assign T_2386 = T_1844 & io_inner_release_bits_voluntary;
  assign T_2392_0 = 4'h0;
  assign T_2392_1 = 4'h8;
  assign T_2394 = T_2392_0 == T_55;
  assign T_2395 = T_2392_1 == T_55;
  assign T_2398 = T_2394 | T_2395;
  assign T_2400 = T_2398 == 1'h0;
  assign T_2401 = T_2386 & T_2400;
  assign T_2403 = T_44 == 1'h0;
  assign T_2404 = T_2401 & T_2403;
  assign T_2405 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2407 = T_2405 == 1'h0;
  assign T_2408 = T_2404 & T_2407;
  assign T_2411 = T_2321 == 1'h0;
  assign T_2412 = T_2408 & T_2411;
  assign T_2414 = T_144_pending == 1'h0;
  assign T_2415 = T_2412 & T_2414;
  assign T_2422_0 = 3'h0;
  assign T_2422_1 = 3'h1;
  assign T_2422_2 = 3'h2;
  assign T_2424 = T_2422_0 == io_inner_release_bits_r_type;
  assign T_2425 = T_2422_1 == io_inner_release_bits_r_type;
  assign T_2426 = T_2422_2 == io_inner_release_bits_r_type;
  assign T_2429 = T_2424 | T_2425;
  assign T_2430 = T_2429 | T_2426;
  assign T_2433 = T_2430 == 1'h0;
  assign T_2435 = io_inner_release_bits_addr_beat == GEN_433;
  assign T_2436 = T_2433 | T_2435;
  assign T_2437 = T_2415 & T_2436;
  assign T_2438 = io_alloc_irel_should | T_2437;
  assign T_2445_0 = 3'h0;
  assign T_2445_1 = 3'h1;
  assign T_2445_2 = 3'h2;
  assign T_2447 = T_2445_0 == io_inner_release_bits_r_type;
  assign T_2448 = T_2445_1 == io_inner_release_bits_r_type;
  assign T_2449 = T_2445_2 == io_inner_release_bits_r_type;
  assign T_2452 = T_2447 | T_2448;
  assign T_2453 = T_2452 | T_2449;
  assign T_2461_0 = 3'h0;
  assign T_2461_1 = 3'h1;
  assign T_2461_2 = 3'h2;
  assign T_2463 = T_2461_0 == io_inner_release_bits_r_type;
  assign T_2464 = T_2461_1 == io_inner_release_bits_r_type;
  assign T_2465 = T_2461_2 == io_inner_release_bits_r_type;
  assign T_2468 = T_2463 | T_2464;
  assign T_2469 = T_2468 | T_2465;
  assign T_2470 = T_2228 & T_2469;
  assign GEN_458 = {{7'd0}, T_2470};
  assign T_2472 = 8'h0 - GEN_458;
  assign T_2473 = T_2472[7:0];
  assign T_2474 = ~ T_2473;
  assign T_2476 = GEN_437 << io_inner_release_bits_addr_beat;
  assign T_2477 = ~ T_2476;
  assign T_2478 = T_2474 | T_2477;
  assign T_2480 = T_2453 ? T_2478 : {{7'd0}, 1'h0};
  assign GEN_56 = T_2438 ? io_inner_release_bits_r_type : T_129;
  assign GEN_57 = T_2438 ? io_inner_release_bits_client_id : T_131;
  assign GEN_58 = T_2438 ? io_inner_release_bits_client_xact_id : T_133;
  assign GEN_65 = T_2438 ? T_2480 : T_135;
  assign T_2484 = T_1844 & T_2231;
  assign T_2486 = T_2484 & T_2208;
  assign T_2488 = T_2438 == 1'h0;
  assign T_2489 = T_2488 & T_2486;
  assign T_2496_0 = 3'h0;
  assign T_2496_1 = 3'h1;
  assign T_2496_2 = 3'h2;
  assign T_2498 = T_2496_0 == io_inner_release_bits_r_type;
  assign T_2499 = T_2496_1 == io_inner_release_bits_r_type;
  assign T_2500 = T_2496_2 == io_inner_release_bits_r_type;
  assign T_2503 = T_2498 | T_2499;
  assign T_2504 = T_2503 | T_2500;
  assign T_2505 = T_2228 & T_2504;
  assign GEN_460 = {{7'd0}, T_2505};
  assign T_2507 = 8'h0 - GEN_460;
  assign T_2508 = T_2507[7:0];
  assign T_2509 = ~ T_2508;
  assign T_2513 = T_2509 | T_2477;
  assign T_2514 = T_135 & T_2513;
  assign GEN_69 = T_2489 ? T_2514 : GEN_65;
  assign GEN_75 = T_2228 ? GEN_56 : T_129;
  assign GEN_76 = T_2228 ? GEN_57 : T_131;
  assign GEN_77 = T_2228 ? GEN_58 : T_133;
  assign GEN_84 = T_2228 ? GEN_69 : T_135;
  assign T_2520_0 = 4'h3;
  assign T_2520_1 = 4'h4;
  assign T_2520_2 = 4'h5;
  assign T_2520_3 = 4'h7;
  assign T_2522 = T_2520_0 == T_55;
  assign T_2523 = T_2520_1 == T_55;
  assign T_2524 = T_2520_2 == T_55;
  assign T_2525 = T_2520_3 == T_55;
  assign T_2528 = T_2522 | T_2523;
  assign T_2529 = T_2528 | T_2524;
  assign T_2530 = T_2529 | T_2525;
  assign T_2531 = T_2530 & T_144_pending;
  assign T_2533 = T_135 != GEN_432;
  assign T_2534 = T_2533 | T_210_pending;
  assign T_2536 = T_2534 == 1'h0;
  assign T_2537 = T_2531 & T_2536;
  assign T_2572_addr_beat = {{2'd0}, 1'h0};
  assign T_2572_addr_block = T_57;
  assign T_2572_client_xact_id = T_133;
  assign T_2572_voluntary = 1'h1;
  assign T_2572_r_type = T_129;
  assign T_2572_data = {{63'd0}, 1'h0};
  assign T_2572_client_id = T_131;
  assign T_2639_addr_beat = {{2'd0}, 1'h0};
  assign T_2639_client_xact_id = T_2572_client_xact_id;
  assign T_2639_manager_xact_id = {{2'd0}, 1'h0};
  assign T_2639_is_builtin_type = 1'h1;
  assign T_2639_g_type = {{1'd0}, 3'h0};
  assign T_2639_data = {{63'd0}, 1'h0};
  assign T_2639_client_id = T_2572_client_id;
  assign T_2679_0 = 4'h0;
  assign T_2679_1 = 4'h8;
  assign T_2681 = T_2679_0 == T_55;
  assign T_2682 = T_2679_1 == T_55;
  assign T_2685 = T_2681 | T_2682;
  assign T_2687 = T_2685 == 1'h0;
  assign T_2688 = T_2386 & T_2687;
  assign T_2691 = T_2688 & T_2403;
  assign T_2695 = T_2691 & T_2407;
  assign T_2699 = T_2695 & T_2411;
  assign T_2702 = T_2699 & T_2414;
  assign T_2709 = T_2702 | T_2486;
  assign T_2716_0 = 3'h0;
  assign T_2716_1 = 3'h1;
  assign T_2716_2 = 3'h2;
  assign T_2718 = T_2716_0 == io_inner_release_bits_r_type;
  assign T_2719 = T_2716_1 == io_inner_release_bits_r_type;
  assign T_2720 = T_2716_2 == io_inner_release_bits_r_type;
  assign T_2723 = T_2718 | T_2719;
  assign T_2724 = T_2723 | T_2720;
  assign T_2725 = T_2228 & T_2724;
  assign GEN_0 = GEN_94;
  assign GEN_88 = GEN_444 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_465 = {{1'd0}, 2'h2};
  assign GEN_89 = GEN_465 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_88;
  assign GEN_466 = {{1'd0}, 2'h3};
  assign GEN_90 = GEN_466 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_89;
  assign GEN_91 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_90;
  assign GEN_92 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_91;
  assign GEN_93 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_92;
  assign GEN_94 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_93;
  assign T_2726 = GEN_0[0];
  assign GEN_1 = GEN_94;
  assign T_2727 = GEN_1[1];
  assign GEN_2 = GEN_94;
  assign T_2728 = GEN_2[2];
  assign GEN_3 = GEN_94;
  assign T_2729 = GEN_3[3];
  assign GEN_4 = GEN_94;
  assign T_2730 = GEN_4[4];
  assign GEN_5 = GEN_94;
  assign T_2731 = GEN_5[5];
  assign GEN_6 = GEN_94;
  assign T_2732 = GEN_6[6];
  assign GEN_7 = GEN_94;
  assign T_2733 = GEN_7[7];
  assign GEN_488 = {{7'd0}, T_2726};
  assign T_2735 = 8'h0 - GEN_488;
  assign T_2736 = T_2735[7:0];
  assign GEN_489 = {{7'd0}, T_2727};
  assign T_2738 = 8'h0 - GEN_489;
  assign T_2739 = T_2738[7:0];
  assign GEN_490 = {{7'd0}, T_2728};
  assign T_2741 = 8'h0 - GEN_490;
  assign T_2742 = T_2741[7:0];
  assign GEN_491 = {{7'd0}, T_2729};
  assign T_2744 = 8'h0 - GEN_491;
  assign T_2745 = T_2744[7:0];
  assign GEN_492 = {{7'd0}, T_2730};
  assign T_2747 = 8'h0 - GEN_492;
  assign T_2748 = T_2747[7:0];
  assign GEN_493 = {{7'd0}, T_2731};
  assign T_2750 = 8'h0 - GEN_493;
  assign T_2751 = T_2750[7:0];
  assign GEN_494 = {{7'd0}, T_2732};
  assign T_2753 = 8'h0 - GEN_494;
  assign T_2754 = T_2753[7:0];
  assign GEN_495 = {{7'd0}, T_2733};
  assign T_2756 = 8'h0 - GEN_495;
  assign T_2757 = T_2756[7:0];
  assign T_2763_0 = T_2736;
  assign T_2763_1 = T_2739;
  assign T_2763_2 = T_2742;
  assign T_2763_3 = T_2745;
  assign T_2763_4 = T_2748;
  assign T_2763_5 = T_2751;
  assign T_2763_6 = T_2754;
  assign T_2763_7 = T_2757;
  assign T_2765 = {T_2763_1,T_2763_0};
  assign T_2766 = {T_2763_3,T_2763_2};
  assign T_2767 = {T_2766,T_2765};
  assign T_2768 = {T_2763_5,T_2763_4};
  assign T_2769 = {T_2763_7,T_2763_6};
  assign T_2770 = {T_2769,T_2768};
  assign T_2771 = {T_2770,T_2767};
  assign T_2772 = ~ T_2771;
  assign T_2773 = T_2772 & io_inner_release_bits_data;
  assign GEN_8 = GEN_150;
  assign GEN_144 = GEN_444 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_145 = GEN_465 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_144;
  assign GEN_146 = GEN_466 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_145;
  assign GEN_147 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_146;
  assign GEN_148 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_147;
  assign GEN_149 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_148;
  assign GEN_150 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_149;
  assign T_2774 = T_2771 & GEN_8;
  assign T_2775 = T_2773 | T_2774;
  assign GEN_9 = T_2775;
  assign GEN_151 = GEN_433 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_152 = GEN_444 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_153 = GEN_465 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_154 = GEN_466 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_155 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_156 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_157 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_158 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_177 = T_2725 ? GEN_151 : data_buffer_0;
  assign GEN_178 = T_2725 ? GEN_152 : data_buffer_1;
  assign GEN_179 = T_2725 ? GEN_153 : data_buffer_2;
  assign GEN_180 = T_2725 ? GEN_154 : data_buffer_3;
  assign GEN_181 = T_2725 ? GEN_155 : data_buffer_4;
  assign GEN_182 = T_2725 ? GEN_156 : data_buffer_5;
  assign GEN_183 = T_2725 ? GEN_157 : data_buffer_6;
  assign GEN_184 = T_2725 ? GEN_158 : data_buffer_7;
  assign T_2806_state = 2'h2;
  assign T_2832 = T_1779 | io_alloc_irel_should;
  assign T_2833 = io_outer_release_ready & io_outer_release_valid;
  assign T_2839_0 = 3'h0;
  assign T_2839_1 = 3'h1;
  assign T_2839_2 = 3'h2;
  assign T_2841 = T_2839_0 == io_outer_release_bits_r_type;
  assign T_2842 = T_2839_1 == io_outer_release_bits_r_type;
  assign T_2843 = T_2839_2 == io_outer_release_bits_r_type;
  assign T_2846 = T_2841 | T_2842;
  assign T_2847 = T_2846 | T_2843;
  assign T_2848 = T_2833 & T_2847;
  assign GEN_503 = {{7'd0}, T_2848};
  assign T_2850 = 8'h0 - GEN_503;
  assign T_2851 = T_2850[7:0];
  assign T_2852 = ~ T_2851;
  assign T_2854 = GEN_437 << io_outer_release_bits_addr_beat;
  assign T_2855 = ~ T_2854;
  assign T_2856 = T_2852 | T_2855;
  assign T_2857 = T_201 & T_2856;
  assign T_2865_0 = 3'h0;
  assign T_2865_1 = 3'h1;
  assign T_2865_2 = 3'h2;
  assign T_2867 = T_2865_0 == io_inner_release_bits_r_type;
  assign T_2868 = T_2865_1 == io_inner_release_bits_r_type;
  assign T_2869 = T_2865_2 == io_inner_release_bits_r_type;
  assign T_2872 = T_2867 | T_2868;
  assign T_2873 = T_2872 | T_2869;
  assign T_2874 = T_2228 & T_2873;
  assign GEN_505 = {{7'd0}, T_2874};
  assign T_2877 = 8'h0 - GEN_505;
  assign T_2878 = T_2877[7:0];
  assign T_2881 = T_2878 & T_2476;
  assign T_2882 = T_2857 | T_2881;
  assign T_2883 = T_2882 | GEN_432;
  assign GEN_191 = T_2832 ? T_2883 : T_201;
  assign GEN_193 = T_2833 ? 1'h0 : T_199;
  assign T_2893 = T_2833 & io_outer_release_bits_voluntary;
  assign T_2900_0 = 3'h0;
  assign T_2900_1 = 3'h1;
  assign T_2900_2 = 3'h2;
  assign T_2902 = T_2900_0 == io_outer_release_bits_r_type;
  assign T_2903 = T_2900_1 == io_outer_release_bits_r_type;
  assign T_2904 = T_2900_2 == io_outer_release_bits_r_type;
  assign T_2907 = T_2902 | T_2903;
  assign T_2908 = T_2907 | T_2904;
  assign T_2910 = T_2893 & T_2908;
  assign T_2914 = T_2912 == 3'h7;
  assign T_2916 = T_2912 + GEN_444;
  assign T_2917 = T_2916[2:0];
  assign GEN_194 = T_2910 ? T_2917 : T_2912;
  assign T_2918 = T_2910 & T_2914;
  assign T_2919 = T_2908 ? T_2912 : {{2'd0}, 1'h0};
  assign T_2920 = T_2908 ? T_2918 : T_2893;
  assign T_2923 = io_outer_grant_bits_g_type == GEN_452;
  assign T_2924 = io_outer_grant_bits_is_builtin_type & T_2923;
  assign T_2925 = T_2405 & T_2924;
  assign T_2933_0 = 3'h5;
  assign GEN_510 = {{1'd0}, T_2933_0};
  assign T_2935 = GEN_510 == io_outer_grant_bits_g_type;
  assign T_2943_0 = 1'h0;
  assign GEN_511 = {{3'd0}, T_2943_0};
  assign T_2945 = GEN_511 == io_outer_grant_bits_g_type;
  assign T_2948 = io_outer_grant_bits_is_builtin_type ? T_2935 : T_2945;
  assign T_2950 = T_2925 & T_2948;
  assign T_2954 = T_2952 == 3'h7;
  assign T_2956 = T_2952 + GEN_444;
  assign T_2957 = T_2956[2:0];
  assign GEN_195 = T_2950 ? T_2957 : T_2952;
  assign T_2958 = T_2950 & T_2954;
  assign T_2959 = T_2948 ? T_2952 : {{2'd0}, 1'h0};
  assign T_2960 = T_2948 ? T_2958 : T_2925;
  assign T_2964 = T_2960 == 1'h0;
  assign T_2965 = T_2920 & T_2964;
  assign T_2967 = T_2962 + 1'h1;
  assign T_2968 = T_2967[0:0];
  assign GEN_196 = T_2965 ? T_2968 : T_2962;
  assign T_2970 = T_2920 == 1'h0;
  assign T_2971 = T_2960 & T_2970;
  assign T_2973 = T_2962 - 1'h1;
  assign T_2974 = T_2973[0:0];
  assign GEN_197 = T_2971 ? T_2974 : GEN_196;
  assign T_2976 = T_2962 > 1'h0;
  assign T_2977 = T_55 == 4'h7;
  assign T_2983_0 = 3'h0;
  assign T_2983_1 = 3'h1;
  assign T_2983_2 = 3'h2;
  assign T_2985 = T_2983_0 == io_outer_release_bits_r_type;
  assign T_2986 = T_2983_1 == io_outer_release_bits_r_type;
  assign T_2987 = T_2983_2 == io_outer_release_bits_r_type;
  assign T_2990 = T_2985 | T_2986;
  assign T_2991 = T_2990 | T_2987;
  assign T_2992 = T_201 >> T_210_up_idx;
  assign T_2993 = T_2992[0];
  assign T_2995 = T_2991 ? T_2993 : T_221;
  assign T_2996 = T_2977 & T_2995;
  assign T_3004_0 = 2'h2;
  assign T_3006 = T_3004_0 == T_2806_state;
  assign T_3009 = T_3006 ? 3'h0 : 3'h3;
  assign T_3045_addr_beat = T_210_up_idx;
  assign T_3045_addr_block = T_57;
  assign T_3045_client_xact_id = {{2'd0}, 1'h0};
  assign T_3045_voluntary = 1'h1;
  assign T_3045_r_type = T_3009;
  assign T_3045_data = GEN_10;
  assign GEN_10 = GEN_204;
  assign GEN_198 = GEN_444 == T_210_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_199 = GEN_465 == T_210_up_idx ? data_buffer_2 : GEN_198;
  assign GEN_200 = GEN_466 == T_210_up_idx ? data_buffer_3 : GEN_199;
  assign GEN_201 = 3'h4 == T_210_up_idx ? data_buffer_4 : GEN_200;
  assign GEN_202 = 3'h5 == T_210_up_idx ? data_buffer_5 : GEN_201;
  assign GEN_203 = 3'h6 == T_210_up_idx ? data_buffer_6 : GEN_202;
  assign GEN_204 = 3'h7 == T_210_up_idx ? data_buffer_7 : GEN_203;
  assign T_3074 = T_99_is_builtin_type == 1'h0;
  assign T_3076 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_3087_0 = 3'h3;
  assign T_3089 = T_3087_0 == io_outer_acquire_bits_a_type;
  assign T_3092 = io_outer_acquire_bits_is_builtin_type & T_3089;
  assign T_3093 = T_3076 & T_3092;
  assign T_3097 = T_3095 == 3'h7;
  assign T_3099 = T_3095 + GEN_444;
  assign T_3100 = T_3099[2:0];
  assign GEN_205 = T_3093 ? T_3100 : T_3095;
  assign T_3101 = T_3093 & T_3097;
  assign T_3102 = T_3092 ? T_3095 : T_69;
  assign T_3103 = T_3092 ? T_3101 : T_3076;
  assign T_3109 = T_2924 == 1'h0;
  assign T_3110 = T_2405 & T_3109;
  assign T_3118_0 = 3'h5;
  assign GEN_518 = {{1'd0}, T_3118_0};
  assign T_3120 = GEN_518 == io_outer_grant_bits_g_type;
  assign T_3128_0 = 1'h0;
  assign GEN_519 = {{3'd0}, T_3128_0};
  assign T_3130 = GEN_519 == io_outer_grant_bits_g_type;
  assign T_3133 = io_outer_grant_bits_is_builtin_type ? T_3120 : T_3130;
  assign T_3135 = T_3110 & T_3133;
  assign T_3139 = T_3137 == 3'h7;
  assign T_3141 = T_3137 + GEN_444;
  assign T_3142 = T_3141[2:0];
  assign GEN_206 = T_3135 ? T_3142 : T_3137;
  assign T_3143 = T_3135 & T_3139;
  assign T_3144 = T_3133 ? T_3137 : T_69;
  assign T_3145 = T_3133 ? T_3143 : T_3110;
  assign T_3149 = T_3145 == 1'h0;
  assign T_3150 = T_3103 & T_3149;
  assign T_3152 = T_3147 + 1'h1;
  assign T_3153 = T_3152[0:0];
  assign GEN_207 = T_3150 ? T_3153 : T_3147;
  assign T_3155 = T_3103 == 1'h0;
  assign T_3156 = T_3145 & T_3155;
  assign T_3158 = T_3147 - 1'h1;
  assign T_3159 = T_3158[0:0];
  assign GEN_208 = T_3156 ? T_3159 : GEN_207;
  assign T_3161 = T_3147 > 1'h0;
  assign T_3162 = T_55 == 4'h6;
  assign T_3163 = T_175 >> T_186_up_idx;
  assign T_3164 = T_3163[0];
  assign T_3166 = T_3164 == 1'h0;
  assign T_3168 = T_59 | T_3166;
  assign T_3169 = T_3162 & T_3168;
  assign T_3172 = T_63 == 5'h1;
  assign T_3173 = T_63 == 5'h7;
  assign T_3174 = T_3172 | T_3173;
  assign T_3175 = T_63[3];
  assign T_3176 = T_63 == 5'h4;
  assign T_3177 = T_3175 | T_3176;
  assign T_3178 = T_3174 | T_3177;
  assign T_3179 = T_63 == 5'h3;
  assign T_3180 = T_3178 | T_3179;
  assign T_3181 = T_63 == 5'h6;
  assign T_3182 = T_3180 | T_3181;
  assign T_3185 = {T_63,1'h1};
  assign T_3216_addr_block = T_57;
  assign T_3216_client_xact_id = {{2'd0}, 1'h0};
  assign T_3216_addr_beat = {{2'd0}, 1'h0};
  assign T_3216_is_builtin_type = 1'h0;
  assign T_3216_a_type = {{2'd0}, T_3182};
  assign T_3216_union = {{6'd0}, T_3185};
  assign T_3216_data = {{63'd0}, 1'h0};
  assign GEN_11 = GEN_215;
  assign GEN_209 = GEN_444 == T_186_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_210 = GEN_465 == T_186_up_idx ? wmask_buffer_2 : GEN_209;
  assign GEN_211 = GEN_466 == T_186_up_idx ? wmask_buffer_3 : GEN_210;
  assign GEN_212 = 3'h4 == T_186_up_idx ? wmask_buffer_4 : GEN_211;
  assign GEN_213 = 3'h5 == T_186_up_idx ? wmask_buffer_5 : GEN_212;
  assign GEN_214 = 3'h6 == T_186_up_idx ? wmask_buffer_6 : GEN_213;
  assign GEN_215 = 3'h7 == T_186_up_idx ? wmask_buffer_7 : GEN_214;
  assign T_3281 = {T_63,1'h0};
  assign T_3282 = {T_65,T_67};
  assign T_3283 = {T_3282,T_3281};
  assign T_3285 = {T_67,T_63};
  assign T_3286 = {T_3285,1'h0};
  assign T_3288 = {GEN_11,1'h0};
  assign T_3300 = T_2111 ? 6'h2 : {{5'd0}, 1'h0};
  assign T_3302 = T_2113 ? 6'h0 : T_3300;
  assign T_3304 = T_2109 ? T_3283 : {{6'd0}, T_3302};
  assign T_3306 = T_2119 ? {{3'd0}, T_3288} : T_3304;
  assign T_3308 = T_2115 ? {{3'd0}, T_3288} : T_3306;
  assign T_3310 = T_2121 ? {{3'd0}, T_3286} : T_3308;
  assign T_3312 = T_2117 ? T_3283 : T_3310;
  assign T_3341_addr_block = T_57;
  assign T_3341_client_xact_id = {{2'd0}, 1'h0};
  assign T_3341_addr_beat = T_186_up_idx;
  assign T_3341_is_builtin_type = 1'h1;
  assign T_3341_a_type = T_99_a_type;
  assign T_3341_union = T_3312;
  assign T_3341_data = GEN_12;
  assign GEN_12 = GEN_222;
  assign GEN_216 = GEN_444 == T_186_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_217 = GEN_465 == T_186_up_idx ? data_buffer_2 : GEN_216;
  assign GEN_218 = GEN_466 == T_186_up_idx ? data_buffer_3 : GEN_217;
  assign GEN_219 = 3'h4 == T_186_up_idx ? data_buffer_4 : GEN_218;
  assign GEN_220 = 3'h5 == T_186_up_idx ? data_buffer_5 : GEN_219;
  assign GEN_221 = 3'h6 == T_186_up_idx ? data_buffer_6 : GEN_220;
  assign GEN_222 = 3'h7 == T_186_up_idx ? data_buffer_7 : GEN_221;
  assign T_3369_addr_block = T_3074 ? T_3216_addr_block : T_3341_addr_block;
  assign T_3369_client_xact_id = T_3074 ? T_3216_client_xact_id : T_3341_client_xact_id;
  assign T_3369_addr_beat = T_3074 ? T_3216_addr_beat : T_3341_addr_beat;
  assign T_3369_is_builtin_type = T_3074 ? T_3216_is_builtin_type : T_3341_is_builtin_type;
  assign T_3369_a_type = T_3074 ? T_3216_a_type : T_3341_a_type;
  assign T_3369_union = T_3074 ? T_3216_union : T_3341_union;
  assign T_3369_data = T_3074 ? T_3216_data : T_3341_data;
  assign T_3398 = T_3162 & T_186_up_done;
  assign GEN_223 = T_3398 ? 4'h7 : GEN_55;
  assign T_3408_0 = 3'h5;
  assign T_3408_1 = 3'h4;
  assign GEN_527 = {{1'd0}, T_3408_0};
  assign T_3410 = GEN_527 == io_outer_grant_bits_g_type;
  assign GEN_528 = {{1'd0}, T_3408_1};
  assign T_3411 = GEN_528 == io_outer_grant_bits_g_type;
  assign T_3414 = T_3410 | T_3411;
  assign T_3420_0 = 1'h0;
  assign GEN_529 = {{3'd0}, T_3420_0};
  assign T_3422 = GEN_529 == io_outer_grant_bits_g_type;
  assign T_3425 = io_outer_grant_bits_is_builtin_type ? T_3414 : T_3422;
  assign T_3426 = T_2405 & T_3425;
  assign GEN_13 = GEN_230;
  assign GEN_224 = GEN_444 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_225 = GEN_465 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_224;
  assign GEN_226 = GEN_466 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_225;
  assign GEN_227 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_226;
  assign GEN_228 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_227;
  assign GEN_229 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_228;
  assign GEN_230 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_229;
  assign T_3427 = GEN_13[0];
  assign GEN_14 = GEN_230;
  assign T_3428 = GEN_14[1];
  assign GEN_15 = GEN_230;
  assign T_3429 = GEN_15[2];
  assign GEN_16 = GEN_230;
  assign T_3430 = GEN_16[3];
  assign GEN_17 = GEN_230;
  assign T_3431 = GEN_17[4];
  assign GEN_18 = GEN_230;
  assign T_3432 = GEN_18[5];
  assign GEN_19 = GEN_230;
  assign T_3433 = GEN_19[6];
  assign GEN_20 = GEN_230;
  assign T_3434 = GEN_20[7];
  assign GEN_554 = {{7'd0}, T_3427};
  assign T_3436 = 8'h0 - GEN_554;
  assign T_3437 = T_3436[7:0];
  assign GEN_555 = {{7'd0}, T_3428};
  assign T_3439 = 8'h0 - GEN_555;
  assign T_3440 = T_3439[7:0];
  assign GEN_556 = {{7'd0}, T_3429};
  assign T_3442 = 8'h0 - GEN_556;
  assign T_3443 = T_3442[7:0];
  assign GEN_557 = {{7'd0}, T_3430};
  assign T_3445 = 8'h0 - GEN_557;
  assign T_3446 = T_3445[7:0];
  assign GEN_558 = {{7'd0}, T_3431};
  assign T_3448 = 8'h0 - GEN_558;
  assign T_3449 = T_3448[7:0];
  assign GEN_559 = {{7'd0}, T_3432};
  assign T_3451 = 8'h0 - GEN_559;
  assign T_3452 = T_3451[7:0];
  assign GEN_560 = {{7'd0}, T_3433};
  assign T_3454 = 8'h0 - GEN_560;
  assign T_3455 = T_3454[7:0];
  assign GEN_561 = {{7'd0}, T_3434};
  assign T_3457 = 8'h0 - GEN_561;
  assign T_3458 = T_3457[7:0];
  assign T_3464_0 = T_3437;
  assign T_3464_1 = T_3440;
  assign T_3464_2 = T_3443;
  assign T_3464_3 = T_3446;
  assign T_3464_4 = T_3449;
  assign T_3464_5 = T_3452;
  assign T_3464_6 = T_3455;
  assign T_3464_7 = T_3458;
  assign T_3466 = {T_3464_1,T_3464_0};
  assign T_3467 = {T_3464_3,T_3464_2};
  assign T_3468 = {T_3467,T_3466};
  assign T_3469 = {T_3464_5,T_3464_4};
  assign T_3470 = {T_3464_7,T_3464_6};
  assign T_3471 = {T_3470,T_3469};
  assign T_3472 = {T_3471,T_3468};
  assign T_3473 = ~ T_3472;
  assign T_3474 = T_3473 & io_outer_grant_bits_data;
  assign GEN_21 = GEN_286;
  assign GEN_280 = GEN_444 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_281 = GEN_465 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_280;
  assign GEN_282 = GEN_466 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_281;
  assign GEN_283 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_282;
  assign GEN_284 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_283;
  assign GEN_285 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_284;
  assign GEN_286 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_285;
  assign T_3475 = T_3472 & GEN_21;
  assign T_3476 = T_3474 | T_3475;
  assign GEN_22 = T_3476;
  assign GEN_287 = GEN_433 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_177;
  assign GEN_288 = GEN_444 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_178;
  assign GEN_289 = GEN_465 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_179;
  assign GEN_290 = GEN_466 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_180;
  assign GEN_291 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_181;
  assign GEN_292 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_182;
  assign GEN_293 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_183;
  assign GEN_294 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_184;
  assign GEN_313 = T_3426 ? GEN_287 : GEN_177;
  assign GEN_314 = T_3426 ? GEN_288 : GEN_178;
  assign GEN_315 = T_3426 ? GEN_289 : GEN_179;
  assign GEN_316 = T_3426 ? GEN_290 : GEN_180;
  assign GEN_317 = T_3426 ? GEN_291 : GEN_181;
  assign GEN_318 = T_3426 ? GEN_292 : GEN_182;
  assign GEN_319 = T_3426 ? GEN_293 : GEN_183;
  assign GEN_320 = T_3426 ? GEN_294 : GEN_184;
  assign T_3477 = T_221 | T_186_pending;
  assign T_3478 = T_3477 | T_210_pending;
  assign T_3489 = T_2325 == 1'h0;
  assign T_3491 = T_2321 & T_3489;
  assign T_3499_0 = 3'h5;
  assign GEN_570 = {{1'd0}, T_3499_0};
  assign T_3501 = GEN_570 == io_inner_grant_bits_g_type;
  assign T_3509_0 = 2'h0;
  assign T_3509_1 = 2'h1;
  assign GEN_571 = {{2'd0}, T_3509_0};
  assign T_3511 = GEN_571 == io_inner_grant_bits_g_type;
  assign GEN_572 = {{2'd0}, T_3509_1};
  assign T_3512 = GEN_572 == io_inner_grant_bits_g_type;
  assign T_3515 = T_3511 | T_3512;
  assign T_3516 = io_inner_grant_bits_is_builtin_type ? T_3501 : T_3515;
  assign T_3518 = T_3491 & T_3516;
  assign T_3522 = T_3520 == 3'h7;
  assign T_3524 = T_3520 + GEN_444;
  assign T_3525 = T_3524[2:0];
  assign GEN_321 = T_3518 ? T_3525 : T_3520;
  assign T_3526 = T_3518 & T_3522;
  assign T_3527 = T_3516 ? T_3520 : {{2'd0}, 1'h0};
  assign T_3528 = T_3516 ? T_3526 : T_3491;
  assign T_3529 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3547 = T_3529 == 1'h0;
  assign T_3548 = T_3528 & T_3547;
  assign T_3550 = T_3545 + 1'h1;
  assign T_3551 = T_3550[0:0];
  assign GEN_323 = T_3548 ? T_3551 : T_3545;
  assign T_3553 = T_3528 == 1'h0;
  assign T_3554 = T_3529 & T_3553;
  assign T_3556 = T_3545 - 1'h1;
  assign T_3557 = T_3556[0:0];
  assign GEN_324 = T_3554 ? T_3557 : GEN_323;
  assign T_3559 = T_3545 > 1'h0;
  assign T_3564 = T_1885 == 1'h0;
  assign T_3573_0 = 3'h5;
  assign T_3573_1 = 3'h4;
  assign GEN_575 = {{1'd0}, T_3573_0};
  assign T_3575 = GEN_575 == io_inner_grant_bits_g_type;
  assign GEN_576 = {{1'd0}, T_3573_1};
  assign T_3576 = GEN_576 == io_inner_grant_bits_g_type;
  assign T_3579 = T_3575 | T_3576;
  assign T_3585_0 = 2'h0;
  assign T_3585_1 = 2'h1;
  assign GEN_577 = {{2'd0}, T_3585_0};
  assign T_3587 = GEN_577 == io_inner_grant_bits_g_type;
  assign GEN_578 = {{2'd0}, T_3585_1};
  assign T_3588 = GEN_578 == io_inner_grant_bits_g_type;
  assign T_3591 = T_3587 | T_3588;
  assign T_3592 = io_inner_grant_bits_is_builtin_type ? T_3579 : T_3591;
  assign T_3593 = T_2321 & T_3592;
  assign GEN_579 = {{7'd0}, T_3593};
  assign T_3595 = 8'h0 - GEN_579;
  assign T_3596 = T_3595[7:0];
  assign T_3597 = ~ T_3596;
  assign T_3599 = GEN_437 << io_inner_grant_bits_addr_beat;
  assign T_3600 = ~ T_3599;
  assign T_3601 = T_3597 | T_3600;
  assign T_3602 = T_177 & T_3601;
  assign T_3610_0 = 3'h0;
  assign T_3610_1 = 3'h1;
  assign T_3610_2 = 3'h2;
  assign T_3612 = T_3610_0 == io_inner_release_bits_r_type;
  assign T_3613 = T_3610_1 == io_inner_release_bits_r_type;
  assign T_3614 = T_3610_2 == io_inner_release_bits_r_type;
  assign T_3617 = T_3612 | T_3613;
  assign T_3618 = T_3617 | T_3614;
  assign T_3619 = T_2228 & T_3618;
  assign GEN_581 = {{7'd0}, T_3619};
  assign T_3622 = 8'h0 - GEN_581;
  assign T_3623 = T_3622[7:0];
  assign T_3626 = T_3623 & T_2476;
  assign T_3627 = T_3602 | T_3626;
  assign T_3637_0 = 3'h5;
  assign T_3637_1 = 3'h4;
  assign GEN_583 = {{1'd0}, T_3637_0};
  assign T_3639 = GEN_583 == io_outer_grant_bits_g_type;
  assign GEN_584 = {{1'd0}, T_3637_1};
  assign T_3640 = GEN_584 == io_outer_grant_bits_g_type;
  assign T_3643 = T_3639 | T_3640;
  assign T_3649_0 = 1'h0;
  assign GEN_585 = {{3'd0}, T_3649_0};
  assign T_3651 = GEN_585 == io_outer_grant_bits_g_type;
  assign T_3654 = io_outer_grant_bits_is_builtin_type ? T_3643 : T_3651;
  assign T_3655 = T_2405 & T_3654;
  assign GEN_586 = {{7'd0}, T_3655};
  assign T_3658 = 8'h0 - GEN_586;
  assign T_3659 = T_3658[7:0];
  assign T_3661 = GEN_437 << io_outer_grant_bits_addr_beat;
  assign T_3662 = T_3659 & T_3661;
  assign T_3663 = T_3627 | T_3662;
  assign T_3664 = T_3663 | GEN_432;
  assign GEN_335 = T_3564 ? T_3664 : GEN_43;
  assign T_3666 = T_55 == 4'h1;
  assign T_3667 = T_1733 | T_3666;
  assign T_3670 = T_3667 | T_2075;
  assign T_3672 = T_3670 == 1'h0;
  assign T_3689 = 3'h6 == Queue_13_1_io_deq_bits_a_type;
  assign T_3690 = T_3689 ? 3'h1 : 3'h3;
  assign T_3691 = 3'h5 == Queue_13_1_io_deq_bits_a_type;
  assign T_3692 = T_3691 ? 3'h1 : T_3690;
  assign T_3693 = 3'h4 == Queue_13_1_io_deq_bits_a_type;
  assign T_3694 = T_3693 ? 3'h4 : T_3692;
  assign T_3695 = 3'h3 == Queue_13_1_io_deq_bits_a_type;
  assign T_3696 = T_3695 ? 3'h3 : T_3694;
  assign T_3697 = 3'h2 == Queue_13_1_io_deq_bits_a_type;
  assign T_3698 = T_3697 ? 3'h3 : T_3696;
  assign T_3699 = 3'h1 == Queue_13_1_io_deq_bits_a_type;
  assign T_3700 = T_3699 ? 3'h5 : T_3698;
  assign T_3701 = 3'h0 == Queue_13_1_io_deq_bits_a_type;
  assign T_3702 = T_3701 ? 3'h4 : T_3700;
  assign T_3703 = Queue_13_1_io_deq_bits_a_type == GEN_433;
  assign T_3708 = T_3703 ? 2'h0 : 2'h1;
  assign T_3709 = Queue_13_1_io_deq_bits_is_builtin_type ? T_3702 : {{1'd0}, T_3708};
  assign T_3741_addr_beat = Queue_13_1_io_deq_bits_addr_beat;
  assign T_3741_client_xact_id = Queue_13_1_io_deq_bits_client_xact_id;
  assign T_3741_manager_xact_id = {{1'd0}, 2'h3};
  assign T_3741_is_builtin_type = Queue_13_1_io_deq_bits_is_builtin_type;
  assign T_3741_g_type = {{1'd0}, T_3709};
  assign T_3741_data = GEN_23;
  assign T_3741_client_id = Queue_13_1_io_deq_bits_client_id;
  assign GEN_23 = GEN_342;
  assign GEN_336 = GEN_444 == T_155 ? data_buffer_1 : data_buffer_0;
  assign GEN_337 = GEN_465 == T_155 ? data_buffer_2 : GEN_336;
  assign GEN_338 = GEN_466 == T_155 ? data_buffer_3 : GEN_337;
  assign GEN_339 = 3'h4 == T_155 ? data_buffer_4 : GEN_338;
  assign GEN_340 = 3'h5 == T_155 ? data_buffer_5 : GEN_339;
  assign GEN_341 = 3'h6 == T_155 ? data_buffer_6 : GEN_340;
  assign GEN_342 = 3'h7 == T_155 ? data_buffer_7 : GEN_341;
  assign T_3780_0 = 3'h5;
  assign GEN_594 = {{1'd0}, T_3780_0};
  assign T_3782 = GEN_594 == io_inner_grant_bits_g_type;
  assign T_3790_0 = 2'h0;
  assign T_3790_1 = 2'h1;
  assign GEN_595 = {{2'd0}, T_3790_0};
  assign T_3792 = GEN_595 == io_inner_grant_bits_g_type;
  assign GEN_596 = {{2'd0}, T_3790_1};
  assign T_3793 = GEN_596 == io_inner_grant_bits_g_type;
  assign T_3796 = T_3792 | T_3793;
  assign T_3797 = io_inner_grant_bits_is_builtin_type ? T_3782 : T_3796;
  assign T_3799 = T_2321 & T_3797;
  assign T_3803 = T_3801 == 3'h7;
  assign T_3805 = T_3801 + GEN_444;
  assign T_3806 = T_3805[2:0];
  assign GEN_343 = T_3799 ? T_3806 : T_3801;
  assign T_3807 = T_3799 & T_3803;
  assign T_3808 = T_3797 ? T_3801 : Queue_13_1_io_deq_bits_addr_beat;
  assign T_3809 = T_3797 ? T_3807 : T_2321;
  assign T_3814 = T_2977 & T_153;
  assign T_3816 = T_3478 == 1'h0;
  assign T_3824_0 = 3'h5;
  assign T_3824_1 = 3'h4;
  assign GEN_598 = {{1'd0}, T_3824_0};
  assign T_3826 = GEN_598 == io_inner_grant_bits_g_type;
  assign GEN_599 = {{1'd0}, T_3824_1};
  assign T_3827 = GEN_599 == io_inner_grant_bits_g_type;
  assign T_3830 = T_3826 | T_3827;
  assign T_3836_0 = 2'h0;
  assign T_3836_1 = 2'h1;
  assign GEN_600 = {{2'd0}, T_3836_0};
  assign T_3838 = GEN_600 == io_inner_grant_bits_g_type;
  assign GEN_601 = {{2'd0}, T_3836_1};
  assign T_3839 = GEN_601 == io_inner_grant_bits_g_type;
  assign T_3842 = T_3838 | T_3839;
  assign T_3843 = io_inner_grant_bits_is_builtin_type ? T_3830 : T_3842;
  assign T_3844 = T_177 >> T_155;
  assign T_3845 = T_3844[0];
  assign T_3846 = T_3843 ? T_3845 : T_3672;
  assign T_3847 = T_3816 & T_3846;
  assign GEN_348 = T_3814 ? T_3847 : T_2537;
  assign GEN_349 = T_2414 ? T_157 : 1'h0;
  assign GEN_350 = T_2414 ? T_155 : T_2639_addr_beat;
  assign GEN_351 = T_2414 ? T_3741_client_xact_id : T_2639_client_xact_id;
  assign GEN_352 = T_2414 ? T_3741_manager_xact_id : T_2639_manager_xact_id;
  assign GEN_353 = T_2414 ? T_3741_is_builtin_type : T_2639_is_builtin_type;
  assign GEN_354 = T_2414 ? T_3741_g_type : T_2639_g_type;
  assign GEN_355 = T_2414 ? T_3741_data : T_2639_data;
  assign GEN_356 = T_2414 ? T_3741_client_id : T_2639_client_id;
  assign GEN_361 = T_2414 ? GEN_348 : T_2537;
  assign T_3854 = ~ io_incoherent_0;
  assign GEN_362 = T_1885 ? {{1'd0}, T_3854} : T_2207;
  assign T_3869_0 = 3'h3;
  assign T_3871 = T_3869_0 == T_99_a_type;
  assign T_3874 = T_99_is_builtin_type & T_3871;
  assign T_3875 = T_1887 & T_3874;
  assign T_3876 = T_3875 & T_153;
  assign T_3879 = T_3876 & T_1905;
  assign T_3881 = T_3879 & io_inner_acquire_valid;
  assign T_3882 = T_1885 | T_3881;
  assign T_3892_0 = 3'h2;
  assign T_3892_1 = 3'h3;
  assign T_3892_2 = 3'h4;
  assign T_3894 = T_3892_0 == io_inner_acquire_bits_a_type;
  assign T_3895 = T_3892_1 == io_inner_acquire_bits_a_type;
  assign T_3896 = T_3892_2 == io_inner_acquire_bits_a_type;
  assign T_3899 = T_3894 | T_3895;
  assign T_3900 = T_3899 | T_3896;
  assign T_3901 = io_inner_acquire_bits_is_builtin_type & T_3900;
  assign T_3902 = T_1734 & T_3901;
  assign T_3903 = T_3902 & T_3882;
  assign T_3905 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3906 = io_inner_acquire_bits_is_builtin_type & T_3905;
  assign T_3910 = 8'h0 - GEN_437;
  assign T_3911 = T_3910[7:0];
  assign T_3917_0 = T_3911;
  assign T_3925 = T_2034 | T_2031;
  assign T_3926 = io_inner_acquire_bits_union[8:1];
  assign T_3928 = T_3925 ? T_3926 : {{7'd0}, 1'h0};
  assign T_3929 = T_3906 ? T_3917_0 : T_3928;
  assign T_3930 = T_3929[0];
  assign T_3931 = T_3929[1];
  assign T_3932 = T_3929[2];
  assign T_3933 = T_3929[3];
  assign T_3934 = T_3929[4];
  assign T_3935 = T_3929[5];
  assign T_3936 = T_3929[6];
  assign T_3937 = T_3929[7];
  assign GEN_603 = {{7'd0}, T_3930};
  assign T_3939 = 8'h0 - GEN_603;
  assign T_3940 = T_3939[7:0];
  assign GEN_604 = {{7'd0}, T_3931};
  assign T_3942 = 8'h0 - GEN_604;
  assign T_3943 = T_3942[7:0];
  assign GEN_605 = {{7'd0}, T_3932};
  assign T_3945 = 8'h0 - GEN_605;
  assign T_3946 = T_3945[7:0];
  assign GEN_606 = {{7'd0}, T_3933};
  assign T_3948 = 8'h0 - GEN_606;
  assign T_3949 = T_3948[7:0];
  assign GEN_607 = {{7'd0}, T_3934};
  assign T_3951 = 8'h0 - GEN_607;
  assign T_3952 = T_3951[7:0];
  assign GEN_608 = {{7'd0}, T_3935};
  assign T_3954 = 8'h0 - GEN_608;
  assign T_3955 = T_3954[7:0];
  assign GEN_609 = {{7'd0}, T_3936};
  assign T_3957 = 8'h0 - GEN_609;
  assign T_3958 = T_3957[7:0];
  assign GEN_610 = {{7'd0}, T_3937};
  assign T_3960 = 8'h0 - GEN_610;
  assign T_3961 = T_3960[7:0];
  assign T_3967_0 = T_3940;
  assign T_3967_1 = T_3943;
  assign T_3967_2 = T_3946;
  assign T_3967_3 = T_3949;
  assign T_3967_4 = T_3952;
  assign T_3967_5 = T_3955;
  assign T_3967_6 = T_3958;
  assign T_3967_7 = T_3961;
  assign T_3969 = {T_3967_1,T_3967_0};
  assign T_3970 = {T_3967_3,T_3967_2};
  assign T_3971 = {T_3970,T_3969};
  assign T_3972 = {T_3967_5,T_3967_4};
  assign T_3973 = {T_3967_7,T_3967_6};
  assign T_3974 = {T_3973,T_3972};
  assign T_3975 = {T_3974,T_3971};
  assign T_3976 = ~ T_3975;
  assign GEN_24 = GEN_369;
  assign GEN_363 = GEN_444 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_364 = GEN_465 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_363;
  assign GEN_365 = GEN_466 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_364;
  assign GEN_366 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_365;
  assign GEN_367 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_366;
  assign GEN_368 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_367;
  assign GEN_369 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_368;
  assign T_3977 = T_3976 & GEN_24;
  assign T_3978 = T_3975 & io_inner_acquire_bits_data;
  assign T_3979 = T_3977 | T_3978;
  assign GEN_25 = T_3979;
  assign GEN_370 = GEN_433 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_313;
  assign GEN_371 = GEN_444 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_314;
  assign GEN_372 = GEN_465 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_315;
  assign GEN_373 = GEN_466 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_316;
  assign GEN_374 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_317;
  assign GEN_375 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_318;
  assign GEN_376 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_319;
  assign GEN_377 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_320;
  assign T_3993_0 = T_3911;
  assign T_4005 = T_3906 ? T_3993_0 : T_3928;
  assign GEN_26 = GEN_384;
  assign GEN_378 = GEN_444 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_379 = GEN_465 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_378;
  assign GEN_380 = GEN_466 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_379;
  assign GEN_381 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_380;
  assign GEN_382 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_381;
  assign GEN_383 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_382;
  assign GEN_384 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_383;
  assign T_4006 = T_4005 | GEN_26;
  assign GEN_27 = T_4006;
  assign GEN_385 = GEN_433 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_0;
  assign GEN_386 = GEN_444 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_1;
  assign GEN_387 = GEN_465 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_2;
  assign GEN_388 = GEN_466 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_3;
  assign GEN_389 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_4;
  assign GEN_390 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_5;
  assign GEN_391 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_6;
  assign GEN_392 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_7;
  assign GEN_404 = T_3903 ? GEN_370 : GEN_313;
  assign GEN_405 = T_3903 ? GEN_371 : GEN_314;
  assign GEN_406 = T_3903 ? GEN_372 : GEN_315;
  assign GEN_407 = T_3903 ? GEN_373 : GEN_316;
  assign GEN_408 = T_3903 ? GEN_374 : GEN_317;
  assign GEN_409 = T_3903 ? GEN_375 : GEN_318;
  assign GEN_410 = T_3903 ? GEN_376 : GEN_319;
  assign GEN_411 = T_3903 ? GEN_377 : GEN_320;
  assign GEN_415 = T_3903 ? GEN_385 : wmask_buffer_0;
  assign GEN_416 = T_3903 ? GEN_386 : wmask_buffer_1;
  assign GEN_417 = T_3903 ? GEN_387 : wmask_buffer_2;
  assign GEN_418 = T_3903 ? GEN_388 : wmask_buffer_3;
  assign GEN_419 = T_3903 ? GEN_389 : wmask_buffer_4;
  assign GEN_420 = T_3903 ? GEN_390 : wmask_buffer_5;
  assign GEN_421 = T_3903 ? GEN_391 : wmask_buffer_6;
  assign GEN_422 = T_3903 ? GEN_392 : wmask_buffer_7;
  assign T_4009 = T_2075 | T_2533;
  assign T_4010 = T_4009 | T_144_pending;
  assign T_4011 = T_4010 | T_221;
  assign T_4012 = T_4011 | T_210_pending;
  assign T_4013 = T_4012 | T_186_pending;
  assign T_4014 = T_4013 | T_153;
  assign T_4015 = T_4014 | T_166_pending;
  assign T_4017 = T_4015 == 1'h0;
  assign T_4019 = T_2977 & T_44;
  assign GEN_423 = T_4019 ? 4'h0 : GEN_223;
  assign GEN_424 = T_4019 ? {{7'd0}, 1'h0} : GEN_415;
  assign GEN_425 = T_4019 ? {{7'd0}, 1'h0} : GEN_416;
  assign GEN_426 = T_4019 ? {{7'd0}, 1'h0} : GEN_417;
  assign GEN_427 = T_4019 ? {{7'd0}, 1'h0} : GEN_418;
  assign GEN_428 = T_4019 ? {{7'd0}, 1'h0} : GEN_419;
  assign GEN_429 = T_4019 ? {{7'd0}, 1'h0} : GEN_420;
  assign GEN_430 = T_4019 ? {{7'd0}, 1'h0} : GEN_421;
  assign GEN_431 = T_4019 ? {{7'd0}, 1'h0} : GEN_422;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_30 = {1{$random}};
  T_55 = GEN_30[3:0];
  GEN_31 = {1{$random}};
  T_57 = GEN_31[25:0];
  GEN_39 = {1{$random}};
  T_59 = GEN_39[0:0];
  GEN_40 = {1{$random}};
  T_61 = GEN_40[4:0];
  GEN_41 = {1{$random}};
  T_63 = GEN_41[4:0];
  GEN_45 = {1{$random}};
  T_65 = GEN_45[2:0];
  GEN_59 = {1{$random}};
  T_67 = GEN_59[2:0];
  GEN_60 = {1{$random}};
  T_129 = GEN_60[2:0];
  GEN_61 = {1{$random}};
  T_131 = GEN_61[0:0];
  GEN_62 = {1{$random}};
  T_133 = GEN_62[1:0];
  GEN_63 = {1{$random}};
  T_135 = GEN_63[7:0];
  GEN_64 = {1{$random}};
  T_175 = GEN_64[7:0];
  GEN_66 = {1{$random}};
  T_177 = GEN_66[7:0];
  GEN_67 = {1{$random}};
  T_195 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  T_199 = GEN_68[0:0];
  GEN_70 = {1{$random}};
  T_201 = GEN_70[7:0];
  GEN_71 = {2{$random}};
  data_buffer_0 = GEN_71[63:0];
  GEN_72 = {2{$random}};
  data_buffer_1 = GEN_72[63:0];
  GEN_73 = {2{$random}};
  data_buffer_2 = GEN_73[63:0];
  GEN_74 = {2{$random}};
  data_buffer_3 = GEN_74[63:0];
  GEN_78 = {2{$random}};
  data_buffer_4 = GEN_78[63:0];
  GEN_79 = {2{$random}};
  data_buffer_5 = GEN_79[63:0];
  GEN_80 = {2{$random}};
  data_buffer_6 = GEN_80[63:0];
  GEN_81 = {2{$random}};
  data_buffer_7 = GEN_81[63:0];
  GEN_82 = {1{$random}};
  wmask_buffer_0 = GEN_82[7:0];
  GEN_83 = {1{$random}};
  wmask_buffer_1 = GEN_83[7:0];
  GEN_85 = {1{$random}};
  wmask_buffer_2 = GEN_85[7:0];
  GEN_86 = {1{$random}};
  wmask_buffer_3 = GEN_86[7:0];
  GEN_87 = {1{$random}};
  wmask_buffer_4 = GEN_87[7:0];
  GEN_95 = {1{$random}};
  wmask_buffer_5 = GEN_95[7:0];
  GEN_96 = {1{$random}};
  wmask_buffer_6 = GEN_96[7:0];
  GEN_97 = {1{$random}};
  wmask_buffer_7 = GEN_97[7:0];
  GEN_98 = {1{$random}};
  T_2219 = GEN_98[2:0];
  GEN_99 = {1{$random}};
  T_2252 = GEN_99[2:0];
  GEN_100 = {1{$random}};
  T_2262 = GEN_100[0:0];
  GEN_101 = {1{$random}};
  T_2312 = GEN_101[2:0];
  GEN_102 = {1{$random}};
  T_2356 = GEN_102[2:0];
  GEN_103 = {1{$random}};
  T_2366 = GEN_103[0:0];
  GEN_104 = {1{$random}};
  T_2912 = GEN_104[2:0];
  GEN_105 = {1{$random}};
  T_2952 = GEN_105[2:0];
  GEN_106 = {1{$random}};
  T_2962 = GEN_106[0:0];
  GEN_107 = {1{$random}};
  T_3095 = GEN_107[2:0];
  GEN_108 = {1{$random}};
  T_3137 = GEN_108[2:0];
  GEN_109 = {1{$random}};
  T_3147 = GEN_109[0:0];
  GEN_110 = {1{$random}};
  T_3520 = GEN_110[2:0];
  GEN_111 = {1{$random}};
  T_3535 = GEN_111[2:0];
  GEN_112 = {1{$random}};
  T_3545 = GEN_112[0:0];
  GEN_113 = {1{$random}};
  T_3801 = GEN_113[2:0];
  GEN_114 = {1{$random}};
  GEN_28 = GEN_114[0:0];
  GEN_115 = {1{$random}};
  GEN_29 = GEN_115[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_55 <= 4'h0;
    end else begin
      if(T_4019) begin
        T_55 <= 4'h0;
      end else begin
        if(T_3398) begin
          T_55 <= 4'h7;
        end else begin
          if(T_2383) begin
            T_55 <= 4'h7;
          end else begin
            if(T_2283) begin
              if(T_2183) begin
                T_55 <= 4'h6;
              end else begin
                T_55 <= 4'h7;
              end
            end else begin
              if(T_1885) begin
                T_55 <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_57 <= 26'h0;
    end else begin
      if(T_2383) begin
        T_57 <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1885) begin
          T_57 <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_59 <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_61 <= T_2028;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        if(T_2035) begin
          T_63 <= 5'h1;
        end else begin
          T_63 <= T_2036;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_65 <= T_2038;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_67 <= T_2039;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_129 <= io_inner_release_bits_r_type;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_131 <= io_inner_release_bits_client_id;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_133 <= io_inner_release_bits_client_xact_id;
        end
      end
    end
    if(reset) begin
      T_135 <= 8'h0;
    end else begin
      if(T_2228) begin
        if(T_2489) begin
          T_135 <= T_2514;
        end else begin
          if(T_2438) begin
            if(T_2453) begin
              T_135 <= T_2478;
            end else begin
              T_135 <= {{7'd0}, 1'h0};
            end
          end
        end
      end
    end
    if(reset) begin
      T_175 <= 8'h0;
    end else begin
      if(T_1885) begin
        if(T_2034) begin
          T_175 <= T_2070;
        end else begin
          T_175 <= {{7'd0}, 1'h0};
        end
      end else begin
        if(T_1962) begin
          T_175 <= T_2020;
        end
      end
    end
    if(reset) begin
      T_177 <= 8'h0;
    end else begin
      if(T_3564) begin
        T_177 <= T_3664;
      end else begin
        if(T_1885) begin
          T_177 <= {{7'd0}, 1'h0};
        end
      end
    end
    if(1'h0) begin
    end else begin
      T_195 <= GEN_362[0];
    end
    if(reset) begin
      T_199 <= 1'h0;
    end else begin
      if(T_2833) begin
        T_199 <= 1'h0;
      end
    end
    if(reset) begin
      T_201 <= 8'h0;
    end else begin
      if(T_2832) begin
        T_201 <= T_2883;
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1817_0;
    end else begin
      if(T_3903) begin
        if(GEN_433 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_433 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_433 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_433 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_433 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_433 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_433 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1817_1;
    end else begin
      if(T_3903) begin
        if(GEN_444 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_444 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_444 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_444 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_444 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_444 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_444 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1817_2;
    end else begin
      if(T_3903) begin
        if(GEN_465 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_465 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_465 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_465 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_465 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_465 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_465 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1817_3;
    end else begin
      if(T_3903) begin
        if(GEN_466 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_466 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_466 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_466 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_466 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_466 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_466 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1817_4;
    end else begin
      if(T_3903) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1817_5;
    end else begin
      if(T_3903) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1817_6;
    end else begin
      if(T_3903) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1817_7;
    end else begin
      if(T_3903) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1835_0;
    end else begin
      if(T_4019) begin
        wmask_buffer_0 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_433 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1835_1;
    end else begin
      if(T_4019) begin
        wmask_buffer_1 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_444 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1835_2;
    end else begin
      if(T_4019) begin
        wmask_buffer_2 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_465 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1835_3;
    end else begin
      if(T_4019) begin
        wmask_buffer_3 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_466 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1835_4;
    end else begin
      if(T_4019) begin
        wmask_buffer_4 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1835_5;
    end else begin
      if(T_4019) begin
        wmask_buffer_5 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1835_6;
    end else begin
      if(T_4019) begin
        wmask_buffer_6 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1835_7;
    end else begin
      if(T_4019) begin
        wmask_buffer_7 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      T_2219 <= 3'h0;
    end
    if(reset) begin
      T_2252 <= 3'h0;
    end else begin
      if(T_2250) begin
        T_2252 <= T_2257;
      end
    end
    if(reset) begin
      T_2262 <= 1'h0;
    end else begin
      if(T_2271) begin
        T_2262 <= T_2274;
      end else begin
        if(T_2265) begin
          T_2262 <= T_2268;
        end
      end
    end
    if(reset) begin
      T_2312 <= 3'h0;
    end else begin
      if(T_2310) begin
        T_2312 <= T_2317;
      end
    end
    if(reset) begin
      T_2356 <= 3'h0;
    end else begin
      if(T_2354) begin
        T_2356 <= T_2361;
      end
    end
    if(reset) begin
      T_2366 <= 1'h0;
    end else begin
      if(T_2375) begin
        T_2366 <= T_2378;
      end else begin
        if(T_2369) begin
          T_2366 <= T_2372;
        end
      end
    end
    if(reset) begin
      T_2912 <= 3'h0;
    end else begin
      if(T_2910) begin
        T_2912 <= T_2917;
      end
    end
    if(reset) begin
      T_2952 <= 3'h0;
    end else begin
      if(T_2950) begin
        T_2952 <= T_2957;
      end
    end
    if(reset) begin
      T_2962 <= 1'h0;
    end else begin
      if(T_2971) begin
        T_2962 <= T_2974;
      end else begin
        if(T_2965) begin
          T_2962 <= T_2968;
        end
      end
    end
    if(reset) begin
      T_3095 <= 3'h0;
    end else begin
      if(T_3093) begin
        T_3095 <= T_3100;
      end
    end
    if(reset) begin
      T_3137 <= 3'h0;
    end else begin
      if(T_3135) begin
        T_3137 <= T_3142;
      end
    end
    if(reset) begin
      T_3147 <= 1'h0;
    end else begin
      if(T_3156) begin
        T_3147 <= T_3159;
      end else begin
        if(T_3150) begin
          T_3147 <= T_3153;
        end
      end
    end
    if(reset) begin
      T_3520 <= 3'h0;
    end else begin
      if(T_3518) begin
        T_3520 <= T_3525;
      end
    end
    if(reset) begin
      T_3535 <= 3'h0;
    end
    if(reset) begin
      T_3545 <= 1'h0;
    end else begin
      if(T_3554) begin
        T_3545 <= T_3557;
      end else begin
        if(T_3548) begin
          T_3545 <= T_3551;
        end
      end
    end
    if(reset) begin
      T_3801 <= 3'h0;
    end else begin
      if(T_3799) begin
        T_3801 <= T_3806;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1778) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:95 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1778) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1778) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1792) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:99 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1792) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1792) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1803) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1803) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1803) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BufferedBroadcastAcquireTracker_3(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should
);
  wire  T_44;
  reg [3:0] T_55;
  reg [31:0] GEN_30;
  reg [25:0] T_57;
  reg [31:0] GEN_31;
  reg  T_59;
  reg [31:0] GEN_39;
  reg [4:0] T_61;
  reg [31:0] GEN_40;
  reg [4:0] T_63;
  reg [31:0] GEN_41;
  reg [2:0] T_65;
  reg [31:0] GEN_45;
  reg [2:0] T_67;
  reg [31:0] GEN_59;
  wire [2:0] T_69;
  wire [1:0] T_99_client_xact_id;
  wire [2:0] T_99_addr_beat;
  wire  T_99_client_id;
  wire  T_99_is_builtin_type;
  wire [2:0] T_99_a_type;
  reg [2:0] T_129;
  reg [31:0] GEN_60;
  reg  T_131;
  reg [31:0] GEN_61;
  reg [1:0] T_133;
  reg [31:0] GEN_62;
  reg [7:0] T_135;
  reg [31:0] GEN_63;
  wire  T_144_pending;
  wire [2:0] T_144_up_idx;
  wire  T_144_up_done;
  wire [2:0] T_144_down_idx;
  wire  T_144_down_done;
  wire  T_153;
  wire [2:0] T_155;
  wire  T_157;
  wire  T_166_pending;
  wire [2:0] T_166_up_idx;
  wire  T_166_up_done;
  wire [2:0] T_166_down_idx;
  wire  T_166_down_done;
  reg [7:0] T_175;
  reg [31:0] GEN_64;
  reg [7:0] T_177;
  reg [31:0] GEN_66;
  wire  T_186_pending;
  wire [2:0] T_186_up_idx;
  wire  T_186_up_done;
  wire [2:0] T_186_down_idx;
  wire  T_186_down_done;
  reg  T_195;
  reg [31:0] GEN_67;
  reg  T_199;
  reg [31:0] GEN_68;
  reg [7:0] T_201;
  reg [31:0] GEN_70;
  wire  T_210_pending;
  wire [2:0] T_210_up_idx;
  wire  T_210_up_done;
  wire [2:0] T_210_down_idx;
  wire  T_210_down_done;
  wire [7:0] GEN_432;
  wire  T_219;
  wire  T_220;
  wire  T_221;
  wire  T_247_sharers;
  wire [1:0] T_299_state;
  wire  T_395_inner_sharers;
  wire [1:0] T_395_outer_state;
  wire  T_1733;
  wire  T_1734;
  wire  T_1735;
  wire  T_1736;
  wire [2:0] T_1745_0;
  wire  T_1747;
  wire  T_1750;
  wire  T_1751;
  wire [2:0] T_1760_0;
  wire  T_1762;
  wire  T_1765;
  wire  T_1767;
  wire [2:0] GEN_433;
  wire  T_1769;
  wire  T_1770;
  wire  T_1772;
  wire  T_1773;
  wire  T_1775;
  wire  T_1776;
  wire  T_1778;
  wire  T_1779;
  wire  T_1780;
  wire  T_1782;
  wire  T_1784;
  wire  T_1785;
  wire  T_1786;
  wire  T_1787;
  wire  T_1789;
  wire  T_1790;
  wire  T_1792;
  wire  T_1796;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [63:0] T_1817_0;
  wire [63:0] T_1817_1;
  wire [63:0] T_1817_2;
  wire [63:0] T_1817_3;
  wire [63:0] T_1817_4;
  wire [63:0] T_1817_5;
  wire [63:0] T_1817_6;
  wire [63:0] T_1817_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_71;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_72;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_73;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_74;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_78;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_79;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_80;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_81;
  wire [7:0] T_1835_0;
  wire [7:0] T_1835_1;
  wire [7:0] T_1835_2;
  wire [7:0] T_1835_3;
  wire [7:0] T_1835_4;
  wire [7:0] T_1835_5;
  wire [7:0] T_1835_6;
  wire [7:0] T_1835_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_82;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_83;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_85;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_86;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_87;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_95;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_96;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_97;
  wire  T_1841;
  wire  T_1842;
  wire  T_1844;
  wire  T_1845;
  wire  T_1847;
  wire  T_1848;
  wire  Queue_14_1_clk;
  wire  Queue_14_1_reset;
  wire  Queue_14_1_io_enq_ready;
  wire  Queue_14_1_io_enq_valid;
  wire [1:0] Queue_14_1_io_enq_bits_client_xact_id;
  wire [2:0] Queue_14_1_io_enq_bits_addr_beat;
  wire  Queue_14_1_io_enq_bits_client_id;
  wire  Queue_14_1_io_enq_bits_is_builtin_type;
  wire [2:0] Queue_14_1_io_enq_bits_a_type;
  wire  Queue_14_1_io_deq_ready;
  wire  Queue_14_1_io_deq_valid;
  wire [1:0] Queue_14_1_io_deq_bits_client_xact_id;
  wire [2:0] Queue_14_1_io_deq_bits_addr_beat;
  wire  Queue_14_1_io_deq_bits_client_id;
  wire  Queue_14_1_io_deq_bits_is_builtin_type;
  wire [2:0] Queue_14_1_io_deq_bits_a_type;
  wire [1:0] Queue_14_1_io_count;
  wire  T_1884;
  wire  T_1885;
  wire  T_1887;
  wire [2:0] T_1896_0;
  wire  T_1898;
  wire  T_1901;
  wire  T_1902;
  wire  T_1903;
  wire [7:0] T_1904;
  wire  T_1905;
  wire  T_1906;
  wire  T_1908;
  wire [2:0] T_1917_0;
  wire  T_1919;
  wire  T_1922;
  wire  T_1924;
  wire  T_1927;
  wire  T_1928;
  wire  T_1929;
  wire [1:0] T_1930_client_xact_id;
  wire [2:0] T_1930_addr_beat;
  wire  T_1930_client_id;
  wire  T_1930_is_builtin_type;
  wire [2:0] T_1930_a_type;
  wire [1:0] GEN_435;
  wire  T_1960;
  wire  T_1962;
  wire [2:0] T_1972_0;
  wire [2:0] T_1972_1;
  wire [2:0] T_1972_2;
  wire  T_1974;
  wire  T_1975;
  wire  T_1976;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire  T_1982;
  wire [7:0] GEN_436;
  wire [8:0] T_1984;
  wire [7:0] T_1985;
  wire [7:0] T_1986;
  wire [7:0] GEN_437;
  wire [7:0] T_1988;
  wire [7:0] T_1989;
  wire [7:0] T_1990;
  wire [7:0] T_1991;
  wire [2:0] T_2001_0;
  wire  T_2003;
  wire  T_2006;
  wire  T_2007;
  wire  T_2010;
  wire [7:0] T_2019;
  wire [7:0] T_2020;
  wire [7:0] GEN_32;
  wire [3:0] GEN_439;
  wire [4:0] T_2028;
  wire  T_2030;
  wire  T_2031;
  wire  T_2033;
  wire  T_2034;
  wire  T_2035;
  wire [4:0] T_2036;
  wire [4:0] T_2037;
  wire [2:0] T_2038;
  wire [2:0] T_2039;
  wire [2:0] T_2052_0;
  wire [2:0] T_2052_1;
  wire [2:0] T_2052_2;
  wire  T_2054;
  wire  T_2055;
  wire  T_2056;
  wire  T_2059;
  wire  T_2060;
  wire  T_2061;
  wire  T_2062;
  wire [7:0] GEN_440;
  wire [8:0] T_2064;
  wire [7:0] T_2065;
  wire [7:0] T_2066;
  wire [7:0] T_2070;
  wire [7:0] T_2072;
  wire [25:0] GEN_33;
  wire  GEN_34;
  wire [4:0] GEN_35;
  wire [4:0] GEN_36;
  wire [2:0] GEN_37;
  wire [2:0] GEN_38;
  wire [7:0] GEN_42;
  wire [7:0] GEN_43;
  wire [3:0] GEN_44;
  wire  T_2075;
  wire [2:0] T_2088_0;
  wire  T_2090;
  wire  T_2093;
  wire  T_2094;
  wire  T_2095;
  wire  T_2098;
  wire  T_2099;
  wire [7:0] T_2100;
  wire  skip_outer_acquire;
  wire  T_2109;
  wire [1:0] T_2110;
  wire  T_2111;
  wire [1:0] T_2112;
  wire  T_2113;
  wire [1:0] T_2114;
  wire  T_2115;
  wire [1:0] T_2116;
  wire  T_2117;
  wire [1:0] T_2118;
  wire  T_2119;
  wire [1:0] T_2120;
  wire  T_2121;
  wire [1:0] T_2122;
  wire [2:0] GEN_444;
  wire  T_2123;
  wire [1:0] T_2124;
  wire  T_2125;
  wire [1:0] T_2126;
  wire [1:0] T_2127;
  wire [25:0] T_2155_addr_block;
  wire [1:0] T_2155_p_type;
  wire  T_2155_client_id;
  wire  T_2183;
  wire [3:0] T_2184;
  wire  T_2193_pending;
  wire [2:0] T_2193_up_idx;
  wire  T_2193_up_done;
  wire [2:0] T_2193_down_idx;
  wire  T_2193_down_done;
  wire  T_2201;
  wire  T_2202;
  wire [1:0] GEN_446;
  wire [1:0] T_2204;
  wire [1:0] T_2205;
  wire [1:0] GEN_447;
  wire [1:0] T_2206;
  wire [1:0] GEN_448;
  wire [1:0] T_2207;
  wire  T_2208;
  wire  T_2211;
  reg [2:0] T_2219;
  reg [31:0] GEN_98;
  wire  T_2228;
  wire  T_2231;
  wire  T_2232;
  wire  T_2233;
  wire [2:0] T_2240_0;
  wire [2:0] T_2240_1;
  wire [2:0] T_2240_2;
  wire  T_2242;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  reg [2:0] T_2252;
  reg [31:0] GEN_99;
  wire  T_2254;
  wire [3:0] T_2256;
  wire [2:0] T_2257;
  wire [2:0] GEN_46;
  wire  T_2258;
  wire [2:0] T_2259;
  wire  T_2260;
  reg  T_2262;
  reg [31:0] GEN_100;
  wire  T_2264;
  wire  T_2265;
  wire [1:0] T_2267;
  wire  T_2268;
  wire  GEN_47;
  wire  T_2270;
  wire  T_2271;
  wire [1:0] T_2273;
  wire  T_2274;
  wire  GEN_48;
  wire  T_2276;
  wire  T_2280;
  wire  T_2282;
  wire  T_2283;
  wire [3:0] GEN_49;
  wire  T_2287;
  wire  T_2288;
  wire  T_2293;
  wire [2:0] T_2300_0;
  wire [2:0] T_2300_1;
  wire [2:0] T_2300_2;
  wire  T_2302;
  wire  T_2303;
  wire  T_2304;
  wire  T_2307;
  wire  T_2308;
  wire  T_2310;
  reg [2:0] T_2312;
  reg [31:0] GEN_101;
  wire  T_2314;
  wire [3:0] T_2316;
  wire [2:0] T_2317;
  wire [2:0] GEN_50;
  wire  T_2318;
  wire [2:0] T_2319;
  wire  T_2320;
  wire  T_2321;
  wire [3:0] GEN_452;
  wire  T_2324;
  wire  T_2325;
  wire  T_2326;
  wire  T_2327;
  wire [2:0] T_2335_0;
  wire [3:0] GEN_453;
  wire  T_2337;
  wire [1:0] T_2345_0;
  wire [1:0] T_2345_1;
  wire [3:0] GEN_454;
  wire  T_2347;
  wire [3:0] GEN_455;
  wire  T_2348;
  wire  T_2351;
  wire  T_2352;
  wire  T_2354;
  reg [2:0] T_2356;
  reg [31:0] GEN_102;
  wire  T_2358;
  wire [3:0] T_2360;
  wire [2:0] T_2361;
  wire [2:0] GEN_51;
  wire  T_2362;
  wire [2:0] T_2363;
  wire  T_2364;
  reg  T_2366;
  reg [31:0] GEN_103;
  wire  T_2368;
  wire  T_2369;
  wire [1:0] T_2371;
  wire  T_2372;
  wire  GEN_52;
  wire  T_2374;
  wire  T_2375;
  wire [1:0] T_2377;
  wire  T_2378;
  wire  GEN_53;
  wire  T_2380;
  wire  T_2382;
  wire  T_2383;
  wire [25:0] GEN_54;
  wire [3:0] GEN_55;
  wire  T_2386;
  wire [3:0] T_2392_0;
  wire [3:0] T_2392_1;
  wire  T_2394;
  wire  T_2395;
  wire  T_2398;
  wire  T_2400;
  wire  T_2401;
  wire  T_2403;
  wire  T_2404;
  wire  T_2405;
  wire  T_2407;
  wire  T_2408;
  wire  T_2411;
  wire  T_2412;
  wire  T_2414;
  wire  T_2415;
  wire [2:0] T_2422_0;
  wire [2:0] T_2422_1;
  wire [2:0] T_2422_2;
  wire  T_2424;
  wire  T_2425;
  wire  T_2426;
  wire  T_2429;
  wire  T_2430;
  wire  T_2433;
  wire  T_2435;
  wire  T_2436;
  wire  T_2437;
  wire  T_2438;
  wire [2:0] T_2445_0;
  wire [2:0] T_2445_1;
  wire [2:0] T_2445_2;
  wire  T_2447;
  wire  T_2448;
  wire  T_2449;
  wire  T_2452;
  wire  T_2453;
  wire [2:0] T_2461_0;
  wire [2:0] T_2461_1;
  wire [2:0] T_2461_2;
  wire  T_2463;
  wire  T_2464;
  wire  T_2465;
  wire  T_2468;
  wire  T_2469;
  wire  T_2470;
  wire [7:0] GEN_458;
  wire [8:0] T_2472;
  wire [7:0] T_2473;
  wire [7:0] T_2474;
  wire [7:0] T_2476;
  wire [7:0] T_2477;
  wire [7:0] T_2478;
  wire [7:0] T_2480;
  wire [2:0] GEN_56;
  wire  GEN_57;
  wire [1:0] GEN_58;
  wire [7:0] GEN_65;
  wire  T_2484;
  wire  T_2486;
  wire  T_2488;
  wire  T_2489;
  wire [2:0] T_2496_0;
  wire [2:0] T_2496_1;
  wire [2:0] T_2496_2;
  wire  T_2498;
  wire  T_2499;
  wire  T_2500;
  wire  T_2503;
  wire  T_2504;
  wire  T_2505;
  wire [7:0] GEN_460;
  wire [8:0] T_2507;
  wire [7:0] T_2508;
  wire [7:0] T_2509;
  wire [7:0] T_2513;
  wire [7:0] T_2514;
  wire [7:0] GEN_69;
  wire [2:0] GEN_75;
  wire  GEN_76;
  wire [1:0] GEN_77;
  wire [7:0] GEN_84;
  wire [3:0] T_2520_0;
  wire [3:0] T_2520_1;
  wire [3:0] T_2520_2;
  wire [3:0] T_2520_3;
  wire  T_2522;
  wire  T_2523;
  wire  T_2524;
  wire  T_2525;
  wire  T_2528;
  wire  T_2529;
  wire  T_2530;
  wire  T_2531;
  wire  T_2533;
  wire  T_2534;
  wire  T_2536;
  wire  T_2537;
  wire [2:0] T_2572_addr_beat;
  wire [25:0] T_2572_addr_block;
  wire [1:0] T_2572_client_xact_id;
  wire  T_2572_voluntary;
  wire [2:0] T_2572_r_type;
  wire [63:0] T_2572_data;
  wire  T_2572_client_id;
  wire [2:0] T_2639_addr_beat;
  wire [1:0] T_2639_client_xact_id;
  wire [2:0] T_2639_manager_xact_id;
  wire  T_2639_is_builtin_type;
  wire [3:0] T_2639_g_type;
  wire [63:0] T_2639_data;
  wire  T_2639_client_id;
  wire [3:0] T_2679_0;
  wire [3:0] T_2679_1;
  wire  T_2681;
  wire  T_2682;
  wire  T_2685;
  wire  T_2687;
  wire  T_2688;
  wire  T_2691;
  wire  T_2695;
  wire  T_2699;
  wire  T_2702;
  wire  T_2709;
  wire [2:0] T_2716_0;
  wire [2:0] T_2716_1;
  wire [2:0] T_2716_2;
  wire  T_2718;
  wire  T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [7:0] GEN_0;
  wire [7:0] GEN_88;
  wire [2:0] GEN_465;
  wire [7:0] GEN_89;
  wire [2:0] GEN_466;
  wire [7:0] GEN_90;
  wire [7:0] GEN_91;
  wire [7:0] GEN_92;
  wire [7:0] GEN_93;
  wire [7:0] GEN_94;
  wire  T_2726;
  wire [7:0] GEN_1;
  wire  T_2727;
  wire [7:0] GEN_2;
  wire  T_2728;
  wire [7:0] GEN_3;
  wire  T_2729;
  wire [7:0] GEN_4;
  wire  T_2730;
  wire [7:0] GEN_5;
  wire  T_2731;
  wire [7:0] GEN_6;
  wire  T_2732;
  wire [7:0] GEN_7;
  wire  T_2733;
  wire [7:0] GEN_488;
  wire [8:0] T_2735;
  wire [7:0] T_2736;
  wire [7:0] GEN_489;
  wire [8:0] T_2738;
  wire [7:0] T_2739;
  wire [7:0] GEN_490;
  wire [8:0] T_2741;
  wire [7:0] T_2742;
  wire [7:0] GEN_491;
  wire [8:0] T_2744;
  wire [7:0] T_2745;
  wire [7:0] GEN_492;
  wire [8:0] T_2747;
  wire [7:0] T_2748;
  wire [7:0] GEN_493;
  wire [8:0] T_2750;
  wire [7:0] T_2751;
  wire [7:0] GEN_494;
  wire [8:0] T_2753;
  wire [7:0] T_2754;
  wire [7:0] GEN_495;
  wire [8:0] T_2756;
  wire [7:0] T_2757;
  wire [7:0] T_2763_0;
  wire [7:0] T_2763_1;
  wire [7:0] T_2763_2;
  wire [7:0] T_2763_3;
  wire [7:0] T_2763_4;
  wire [7:0] T_2763_5;
  wire [7:0] T_2763_6;
  wire [7:0] T_2763_7;
  wire [15:0] T_2765;
  wire [15:0] T_2766;
  wire [31:0] T_2767;
  wire [15:0] T_2768;
  wire [15:0] T_2769;
  wire [31:0] T_2770;
  wire [63:0] T_2771;
  wire [63:0] T_2772;
  wire [63:0] T_2773;
  wire [63:0] GEN_8;
  wire [63:0] GEN_144;
  wire [63:0] GEN_145;
  wire [63:0] GEN_146;
  wire [63:0] GEN_147;
  wire [63:0] GEN_148;
  wire [63:0] GEN_149;
  wire [63:0] GEN_150;
  wire [63:0] T_2774;
  wire [63:0] T_2775;
  wire [63:0] GEN_9;
  wire [63:0] GEN_151;
  wire [63:0] GEN_152;
  wire [63:0] GEN_153;
  wire [63:0] GEN_154;
  wire [63:0] GEN_155;
  wire [63:0] GEN_156;
  wire [63:0] GEN_157;
  wire [63:0] GEN_158;
  wire [63:0] GEN_177;
  wire [63:0] GEN_178;
  wire [63:0] GEN_179;
  wire [63:0] GEN_180;
  wire [63:0] GEN_181;
  wire [63:0] GEN_182;
  wire [63:0] GEN_183;
  wire [63:0] GEN_184;
  wire [1:0] T_2806_state;
  wire  T_2832;
  wire  T_2833;
  wire [2:0] T_2839_0;
  wire [2:0] T_2839_1;
  wire [2:0] T_2839_2;
  wire  T_2841;
  wire  T_2842;
  wire  T_2843;
  wire  T_2846;
  wire  T_2847;
  wire  T_2848;
  wire [7:0] GEN_503;
  wire [8:0] T_2850;
  wire [7:0] T_2851;
  wire [7:0] T_2852;
  wire [7:0] T_2854;
  wire [7:0] T_2855;
  wire [7:0] T_2856;
  wire [7:0] T_2857;
  wire [2:0] T_2865_0;
  wire [2:0] T_2865_1;
  wire [2:0] T_2865_2;
  wire  T_2867;
  wire  T_2868;
  wire  T_2869;
  wire  T_2872;
  wire  T_2873;
  wire  T_2874;
  wire [7:0] GEN_505;
  wire [8:0] T_2877;
  wire [7:0] T_2878;
  wire [7:0] T_2881;
  wire [7:0] T_2882;
  wire [7:0] T_2883;
  wire [7:0] GEN_191;
  wire  GEN_193;
  wire  T_2893;
  wire [2:0] T_2900_0;
  wire [2:0] T_2900_1;
  wire [2:0] T_2900_2;
  wire  T_2902;
  wire  T_2903;
  wire  T_2904;
  wire  T_2907;
  wire  T_2908;
  wire  T_2910;
  reg [2:0] T_2912;
  reg [31:0] GEN_104;
  wire  T_2914;
  wire [3:0] T_2916;
  wire [2:0] T_2917;
  wire [2:0] GEN_194;
  wire  T_2918;
  wire [2:0] T_2919;
  wire  T_2920;
  wire  T_2923;
  wire  T_2924;
  wire  T_2925;
  wire [2:0] T_2933_0;
  wire [3:0] GEN_510;
  wire  T_2935;
  wire  T_2943_0;
  wire [3:0] GEN_511;
  wire  T_2945;
  wire  T_2948;
  wire  T_2950;
  reg [2:0] T_2952;
  reg [31:0] GEN_105;
  wire  T_2954;
  wire [3:0] T_2956;
  wire [2:0] T_2957;
  wire [2:0] GEN_195;
  wire  T_2958;
  wire [2:0] T_2959;
  wire  T_2960;
  reg  T_2962;
  reg [31:0] GEN_106;
  wire  T_2964;
  wire  T_2965;
  wire [1:0] T_2967;
  wire  T_2968;
  wire  GEN_196;
  wire  T_2970;
  wire  T_2971;
  wire [1:0] T_2973;
  wire  T_2974;
  wire  GEN_197;
  wire  T_2976;
  wire  T_2977;
  wire [2:0] T_2983_0;
  wire [2:0] T_2983_1;
  wire [2:0] T_2983_2;
  wire  T_2985;
  wire  T_2986;
  wire  T_2987;
  wire  T_2990;
  wire  T_2991;
  wire [7:0] T_2992;
  wire  T_2993;
  wire  T_2995;
  wire  T_2996;
  wire [1:0] T_3004_0;
  wire  T_3006;
  wire [2:0] T_3009;
  wire [2:0] T_3045_addr_beat;
  wire [25:0] T_3045_addr_block;
  wire [2:0] T_3045_client_xact_id;
  wire  T_3045_voluntary;
  wire [2:0] T_3045_r_type;
  wire [63:0] T_3045_data;
  wire [63:0] GEN_10;
  wire [63:0] GEN_198;
  wire [63:0] GEN_199;
  wire [63:0] GEN_200;
  wire [63:0] GEN_201;
  wire [63:0] GEN_202;
  wire [63:0] GEN_203;
  wire [63:0] GEN_204;
  wire  T_3074;
  wire  T_3076;
  wire [2:0] T_3087_0;
  wire  T_3089;
  wire  T_3092;
  wire  T_3093;
  reg [2:0] T_3095;
  reg [31:0] GEN_107;
  wire  T_3097;
  wire [3:0] T_3099;
  wire [2:0] T_3100;
  wire [2:0] GEN_205;
  wire  T_3101;
  wire [2:0] T_3102;
  wire  T_3103;
  wire  T_3109;
  wire  T_3110;
  wire [2:0] T_3118_0;
  wire [3:0] GEN_518;
  wire  T_3120;
  wire  T_3128_0;
  wire [3:0] GEN_519;
  wire  T_3130;
  wire  T_3133;
  wire  T_3135;
  reg [2:0] T_3137;
  reg [31:0] GEN_108;
  wire  T_3139;
  wire [3:0] T_3141;
  wire [2:0] T_3142;
  wire [2:0] GEN_206;
  wire  T_3143;
  wire [2:0] T_3144;
  wire  T_3145;
  reg  T_3147;
  reg [31:0] GEN_109;
  wire  T_3149;
  wire  T_3150;
  wire [1:0] T_3152;
  wire  T_3153;
  wire  GEN_207;
  wire  T_3155;
  wire  T_3156;
  wire [1:0] T_3158;
  wire  T_3159;
  wire  GEN_208;
  wire  T_3161;
  wire  T_3162;
  wire [7:0] T_3163;
  wire  T_3164;
  wire  T_3166;
  wire  T_3168;
  wire  T_3169;
  wire  T_3172;
  wire  T_3173;
  wire  T_3174;
  wire  T_3175;
  wire  T_3176;
  wire  T_3177;
  wire  T_3178;
  wire  T_3179;
  wire  T_3180;
  wire  T_3181;
  wire  T_3182;
  wire [5:0] T_3185;
  wire [25:0] T_3216_addr_block;
  wire [2:0] T_3216_client_xact_id;
  wire [2:0] T_3216_addr_beat;
  wire  T_3216_is_builtin_type;
  wire [2:0] T_3216_a_type;
  wire [11:0] T_3216_union;
  wire [63:0] T_3216_data;
  wire [7:0] GEN_11;
  wire [7:0] GEN_209;
  wire [7:0] GEN_210;
  wire [7:0] GEN_211;
  wire [7:0] GEN_212;
  wire [7:0] GEN_213;
  wire [7:0] GEN_214;
  wire [7:0] GEN_215;
  wire [5:0] T_3281;
  wire [5:0] T_3282;
  wire [11:0] T_3283;
  wire [7:0] T_3285;
  wire [8:0] T_3286;
  wire [8:0] T_3288;
  wire [5:0] T_3300;
  wire [5:0] T_3302;
  wire [11:0] T_3304;
  wire [11:0] T_3306;
  wire [11:0] T_3308;
  wire [11:0] T_3310;
  wire [11:0] T_3312;
  wire [25:0] T_3341_addr_block;
  wire [2:0] T_3341_client_xact_id;
  wire [2:0] T_3341_addr_beat;
  wire  T_3341_is_builtin_type;
  wire [2:0] T_3341_a_type;
  wire [11:0] T_3341_union;
  wire [63:0] T_3341_data;
  wire [63:0] GEN_12;
  wire [63:0] GEN_216;
  wire [63:0] GEN_217;
  wire [63:0] GEN_218;
  wire [63:0] GEN_219;
  wire [63:0] GEN_220;
  wire [63:0] GEN_221;
  wire [63:0] GEN_222;
  wire [25:0] T_3369_addr_block;
  wire [2:0] T_3369_client_xact_id;
  wire [2:0] T_3369_addr_beat;
  wire  T_3369_is_builtin_type;
  wire [2:0] T_3369_a_type;
  wire [11:0] T_3369_union;
  wire [63:0] T_3369_data;
  wire  T_3398;
  wire [3:0] GEN_223;
  wire [2:0] T_3408_0;
  wire [2:0] T_3408_1;
  wire [3:0] GEN_527;
  wire  T_3410;
  wire [3:0] GEN_528;
  wire  T_3411;
  wire  T_3414;
  wire  T_3420_0;
  wire [3:0] GEN_529;
  wire  T_3422;
  wire  T_3425;
  wire  T_3426;
  wire [7:0] GEN_13;
  wire [7:0] GEN_224;
  wire [7:0] GEN_225;
  wire [7:0] GEN_226;
  wire [7:0] GEN_227;
  wire [7:0] GEN_228;
  wire [7:0] GEN_229;
  wire [7:0] GEN_230;
  wire  T_3427;
  wire [7:0] GEN_14;
  wire  T_3428;
  wire [7:0] GEN_15;
  wire  T_3429;
  wire [7:0] GEN_16;
  wire  T_3430;
  wire [7:0] GEN_17;
  wire  T_3431;
  wire [7:0] GEN_18;
  wire  T_3432;
  wire [7:0] GEN_19;
  wire  T_3433;
  wire [7:0] GEN_20;
  wire  T_3434;
  wire [7:0] GEN_554;
  wire [8:0] T_3436;
  wire [7:0] T_3437;
  wire [7:0] GEN_555;
  wire [8:0] T_3439;
  wire [7:0] T_3440;
  wire [7:0] GEN_556;
  wire [8:0] T_3442;
  wire [7:0] T_3443;
  wire [7:0] GEN_557;
  wire [8:0] T_3445;
  wire [7:0] T_3446;
  wire [7:0] GEN_558;
  wire [8:0] T_3448;
  wire [7:0] T_3449;
  wire [7:0] GEN_559;
  wire [8:0] T_3451;
  wire [7:0] T_3452;
  wire [7:0] GEN_560;
  wire [8:0] T_3454;
  wire [7:0] T_3455;
  wire [7:0] GEN_561;
  wire [8:0] T_3457;
  wire [7:0] T_3458;
  wire [7:0] T_3464_0;
  wire [7:0] T_3464_1;
  wire [7:0] T_3464_2;
  wire [7:0] T_3464_3;
  wire [7:0] T_3464_4;
  wire [7:0] T_3464_5;
  wire [7:0] T_3464_6;
  wire [7:0] T_3464_7;
  wire [15:0] T_3466;
  wire [15:0] T_3467;
  wire [31:0] T_3468;
  wire [15:0] T_3469;
  wire [15:0] T_3470;
  wire [31:0] T_3471;
  wire [63:0] T_3472;
  wire [63:0] T_3473;
  wire [63:0] T_3474;
  wire [63:0] GEN_21;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [63:0] GEN_286;
  wire [63:0] T_3475;
  wire [63:0] T_3476;
  wire [63:0] GEN_22;
  wire [63:0] GEN_287;
  wire [63:0] GEN_288;
  wire [63:0] GEN_289;
  wire [63:0] GEN_290;
  wire [63:0] GEN_291;
  wire [63:0] GEN_292;
  wire [63:0] GEN_293;
  wire [63:0] GEN_294;
  wire [63:0] GEN_313;
  wire [63:0] GEN_314;
  wire [63:0] GEN_315;
  wire [63:0] GEN_316;
  wire [63:0] GEN_317;
  wire [63:0] GEN_318;
  wire [63:0] GEN_319;
  wire [63:0] GEN_320;
  wire  T_3477;
  wire  T_3478;
  wire  T_3489;
  wire  T_3491;
  wire [2:0] T_3499_0;
  wire [3:0] GEN_570;
  wire  T_3501;
  wire [1:0] T_3509_0;
  wire [1:0] T_3509_1;
  wire [3:0] GEN_571;
  wire  T_3511;
  wire [3:0] GEN_572;
  wire  T_3512;
  wire  T_3515;
  wire  T_3516;
  wire  T_3518;
  reg [2:0] T_3520;
  reg [31:0] GEN_110;
  wire  T_3522;
  wire [3:0] T_3524;
  wire [2:0] T_3525;
  wire [2:0] GEN_321;
  wire  T_3526;
  wire [2:0] T_3527;
  wire  T_3528;
  wire  T_3529;
  reg [2:0] T_3535;
  reg [31:0] GEN_111;
  reg  T_3545;
  reg [31:0] GEN_112;
  wire  T_3547;
  wire  T_3548;
  wire [1:0] T_3550;
  wire  T_3551;
  wire  GEN_323;
  wire  T_3553;
  wire  T_3554;
  wire [1:0] T_3556;
  wire  T_3557;
  wire  GEN_324;
  wire  T_3559;
  wire  T_3564;
  wire [2:0] T_3573_0;
  wire [2:0] T_3573_1;
  wire [3:0] GEN_575;
  wire  T_3575;
  wire [3:0] GEN_576;
  wire  T_3576;
  wire  T_3579;
  wire [1:0] T_3585_0;
  wire [1:0] T_3585_1;
  wire [3:0] GEN_577;
  wire  T_3587;
  wire [3:0] GEN_578;
  wire  T_3588;
  wire  T_3591;
  wire  T_3592;
  wire  T_3593;
  wire [7:0] GEN_579;
  wire [8:0] T_3595;
  wire [7:0] T_3596;
  wire [7:0] T_3597;
  wire [7:0] T_3599;
  wire [7:0] T_3600;
  wire [7:0] T_3601;
  wire [7:0] T_3602;
  wire [2:0] T_3610_0;
  wire [2:0] T_3610_1;
  wire [2:0] T_3610_2;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3617;
  wire  T_3618;
  wire  T_3619;
  wire [7:0] GEN_581;
  wire [8:0] T_3622;
  wire [7:0] T_3623;
  wire [7:0] T_3626;
  wire [7:0] T_3627;
  wire [2:0] T_3637_0;
  wire [2:0] T_3637_1;
  wire [3:0] GEN_583;
  wire  T_3639;
  wire [3:0] GEN_584;
  wire  T_3640;
  wire  T_3643;
  wire  T_3649_0;
  wire [3:0] GEN_585;
  wire  T_3651;
  wire  T_3654;
  wire  T_3655;
  wire [7:0] GEN_586;
  wire [8:0] T_3658;
  wire [7:0] T_3659;
  wire [7:0] T_3661;
  wire [7:0] T_3662;
  wire [7:0] T_3663;
  wire [7:0] T_3664;
  wire [7:0] GEN_335;
  wire  T_3666;
  wire  T_3667;
  wire  T_3670;
  wire  T_3672;
  wire  T_3689;
  wire [2:0] T_3690;
  wire  T_3691;
  wire [2:0] T_3692;
  wire  T_3693;
  wire [2:0] T_3694;
  wire  T_3695;
  wire [2:0] T_3696;
  wire  T_3697;
  wire [2:0] T_3698;
  wire  T_3699;
  wire [2:0] T_3700;
  wire  T_3701;
  wire [2:0] T_3702;
  wire  T_3703;
  wire [1:0] T_3708;
  wire [2:0] T_3709;
  wire [2:0] T_3741_addr_beat;
  wire [1:0] T_3741_client_xact_id;
  wire [2:0] T_3741_manager_xact_id;
  wire  T_3741_is_builtin_type;
  wire [3:0] T_3741_g_type;
  wire [63:0] T_3741_data;
  wire  T_3741_client_id;
  wire [63:0] GEN_23;
  wire [63:0] GEN_336;
  wire [63:0] GEN_337;
  wire [63:0] GEN_338;
  wire [63:0] GEN_339;
  wire [63:0] GEN_340;
  wire [63:0] GEN_341;
  wire [63:0] GEN_342;
  wire [2:0] T_3780_0;
  wire [3:0] GEN_594;
  wire  T_3782;
  wire [1:0] T_3790_0;
  wire [1:0] T_3790_1;
  wire [3:0] GEN_595;
  wire  T_3792;
  wire [3:0] GEN_596;
  wire  T_3793;
  wire  T_3796;
  wire  T_3797;
  wire  T_3799;
  reg [2:0] T_3801;
  reg [31:0] GEN_113;
  wire  T_3803;
  wire [3:0] T_3805;
  wire [2:0] T_3806;
  wire [2:0] GEN_343;
  wire  T_3807;
  wire [2:0] T_3808;
  wire  T_3809;
  wire  T_3814;
  wire  T_3816;
  wire [2:0] T_3824_0;
  wire [2:0] T_3824_1;
  wire [3:0] GEN_598;
  wire  T_3826;
  wire [3:0] GEN_599;
  wire  T_3827;
  wire  T_3830;
  wire [1:0] T_3836_0;
  wire [1:0] T_3836_1;
  wire [3:0] GEN_600;
  wire  T_3838;
  wire [3:0] GEN_601;
  wire  T_3839;
  wire  T_3842;
  wire  T_3843;
  wire [7:0] T_3844;
  wire  T_3845;
  wire  T_3846;
  wire  T_3847;
  wire  GEN_348;
  wire  GEN_349;
  wire [2:0] GEN_350;
  wire [1:0] GEN_351;
  wire [2:0] GEN_352;
  wire  GEN_353;
  wire [3:0] GEN_354;
  wire [63:0] GEN_355;
  wire  GEN_356;
  wire  GEN_361;
  wire  T_3854;
  wire [1:0] GEN_362;
  wire [2:0] T_3869_0;
  wire  T_3871;
  wire  T_3874;
  wire  T_3875;
  wire  T_3876;
  wire  T_3879;
  wire  T_3881;
  wire  T_3882;
  wire [2:0] T_3892_0;
  wire [2:0] T_3892_1;
  wire [2:0] T_3892_2;
  wire  T_3894;
  wire  T_3895;
  wire  T_3896;
  wire  T_3899;
  wire  T_3900;
  wire  T_3901;
  wire  T_3902;
  wire  T_3903;
  wire  T_3905;
  wire  T_3906;
  wire [8:0] T_3910;
  wire [7:0] T_3911;
  wire [7:0] T_3917_0;
  wire  T_3925;
  wire [7:0] T_3926;
  wire [7:0] T_3928;
  wire [7:0] T_3929;
  wire  T_3930;
  wire  T_3931;
  wire  T_3932;
  wire  T_3933;
  wire  T_3934;
  wire  T_3935;
  wire  T_3936;
  wire  T_3937;
  wire [7:0] GEN_603;
  wire [8:0] T_3939;
  wire [7:0] T_3940;
  wire [7:0] GEN_604;
  wire [8:0] T_3942;
  wire [7:0] T_3943;
  wire [7:0] GEN_605;
  wire [8:0] T_3945;
  wire [7:0] T_3946;
  wire [7:0] GEN_606;
  wire [8:0] T_3948;
  wire [7:0] T_3949;
  wire [7:0] GEN_607;
  wire [8:0] T_3951;
  wire [7:0] T_3952;
  wire [7:0] GEN_608;
  wire [8:0] T_3954;
  wire [7:0] T_3955;
  wire [7:0] GEN_609;
  wire [8:0] T_3957;
  wire [7:0] T_3958;
  wire [7:0] GEN_610;
  wire [8:0] T_3960;
  wire [7:0] T_3961;
  wire [7:0] T_3967_0;
  wire [7:0] T_3967_1;
  wire [7:0] T_3967_2;
  wire [7:0] T_3967_3;
  wire [7:0] T_3967_4;
  wire [7:0] T_3967_5;
  wire [7:0] T_3967_6;
  wire [7:0] T_3967_7;
  wire [15:0] T_3969;
  wire [15:0] T_3970;
  wire [31:0] T_3971;
  wire [15:0] T_3972;
  wire [15:0] T_3973;
  wire [31:0] T_3974;
  wire [63:0] T_3975;
  wire [63:0] T_3976;
  wire [63:0] GEN_24;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [63:0] GEN_366;
  wire [63:0] GEN_367;
  wire [63:0] GEN_368;
  wire [63:0] GEN_369;
  wire [63:0] T_3977;
  wire [63:0] T_3978;
  wire [63:0] T_3979;
  wire [63:0] GEN_25;
  wire [63:0] GEN_370;
  wire [63:0] GEN_371;
  wire [63:0] GEN_372;
  wire [63:0] GEN_373;
  wire [63:0] GEN_374;
  wire [63:0] GEN_375;
  wire [63:0] GEN_376;
  wire [63:0] GEN_377;
  wire [7:0] T_3993_0;
  wire [7:0] T_4005;
  wire [7:0] GEN_26;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [7:0] GEN_381;
  wire [7:0] GEN_382;
  wire [7:0] GEN_383;
  wire [7:0] GEN_384;
  wire [7:0] T_4006;
  wire [7:0] GEN_27;
  wire [7:0] GEN_385;
  wire [7:0] GEN_386;
  wire [7:0] GEN_387;
  wire [7:0] GEN_388;
  wire [7:0] GEN_389;
  wire [7:0] GEN_390;
  wire [7:0] GEN_391;
  wire [7:0] GEN_392;
  wire [63:0] GEN_404;
  wire [63:0] GEN_405;
  wire [63:0] GEN_406;
  wire [63:0] GEN_407;
  wire [63:0] GEN_408;
  wire [63:0] GEN_409;
  wire [63:0] GEN_410;
  wire [63:0] GEN_411;
  wire [7:0] GEN_415;
  wire [7:0] GEN_416;
  wire [7:0] GEN_417;
  wire [7:0] GEN_418;
  wire [7:0] GEN_419;
  wire [7:0] GEN_420;
  wire [7:0] GEN_421;
  wire [7:0] GEN_422;
  wire  T_4009;
  wire  T_4010;
  wire  T_4011;
  wire  T_4012;
  wire  T_4013;
  wire  T_4014;
  wire  T_4015;
  wire  T_4017;
  wire  T_4019;
  wire [3:0] GEN_423;
  wire [7:0] GEN_424;
  wire [7:0] GEN_425;
  wire [7:0] GEN_426;
  wire [7:0] GEN_427;
  wire [7:0] GEN_428;
  wire [7:0] GEN_429;
  wire [7:0] GEN_430;
  wire [7:0] GEN_431;
  reg  GEN_28;
  reg [31:0] GEN_114;
  reg  GEN_29;
  reg [31:0] GEN_115;
  Queue_11 Queue_14_1 (
    .clk(Queue_14_1_clk),
    .reset(Queue_14_1_reset),
    .io_enq_ready(Queue_14_1_io_enq_ready),
    .io_enq_valid(Queue_14_1_io_enq_valid),
    .io_enq_bits_client_xact_id(Queue_14_1_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(Queue_14_1_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(Queue_14_1_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(Queue_14_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(Queue_14_1_io_enq_bits_a_type),
    .io_deq_ready(Queue_14_1_io_deq_ready),
    .io_deq_valid(Queue_14_1_io_deq_valid),
    .io_deq_bits_client_xact_id(Queue_14_1_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(Queue_14_1_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(Queue_14_1_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(Queue_14_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(Queue_14_1_io_deq_bits_a_type),
    .io_count(Queue_14_1_io_count)
  );
  assign io_inner_acquire_ready = T_2099;
  assign io_inner_grant_valid = GEN_361;
  assign io_inner_grant_bits_addr_beat = GEN_350;
  assign io_inner_grant_bits_client_xact_id = GEN_351;
  assign io_inner_grant_bits_manager_xact_id = GEN_352;
  assign io_inner_grant_bits_is_builtin_type = GEN_353;
  assign io_inner_grant_bits_g_type = GEN_354;
  assign io_inner_grant_bits_data = GEN_355;
  assign io_inner_grant_bits_client_id = GEN_356;
  assign io_inner_finish_ready = T_2977;
  assign io_inner_probe_valid = T_2211;
  assign io_inner_probe_bits_addr_block = T_2155_addr_block;
  assign io_inner_probe_bits_p_type = T_2155_p_type;
  assign io_inner_probe_bits_client_id = T_2155_client_id;
  assign io_inner_release_ready = T_2709;
  assign io_outer_acquire_valid = T_3169;
  assign io_outer_acquire_bits_addr_block = T_3369_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3369_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3369_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3369_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3369_a_type;
  assign io_outer_acquire_bits_union = T_3369_union;
  assign io_outer_acquire_bits_data = T_3369_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2996;
  assign io_outer_release_bits_addr_beat = T_3045_addr_beat;
  assign io_outer_release_bits_addr_block = T_3045_addr_block;
  assign io_outer_release_bits_client_xact_id = T_3045_client_xact_id;
  assign io_outer_release_bits_voluntary = T_3045_voluntary;
  assign io_outer_release_bits_r_type = T_3045_r_type;
  assign io_outer_release_bits_data = T_3045_data;
  assign io_outer_grant_ready = T_2977;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_28;
  assign io_outer_finish_bits_manager_id = GEN_29;
  assign io_alloc_iacq_matches = T_1842;
  assign io_alloc_iacq_can = T_1733;
  assign io_alloc_irel_matches = T_1845;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1848;
  assign io_alloc_oprb_can = 1'h0;
  assign T_44 = T_4017;
  assign T_69 = T_99_addr_beat;
  assign T_99_client_xact_id = T_1930_client_xact_id;
  assign T_99_addr_beat = T_1930_addr_beat;
  assign T_99_client_id = T_1930_client_id;
  assign T_99_is_builtin_type = T_1930_is_builtin_type;
  assign T_99_a_type = T_1930_a_type;
  assign T_144_pending = T_2380;
  assign T_144_up_idx = T_2319;
  assign T_144_up_done = T_2320;
  assign T_144_down_idx = T_2363;
  assign T_144_down_done = T_2364;
  assign T_153 = T_1960;
  assign T_155 = T_3808;
  assign T_157 = T_3809;
  assign T_166_pending = T_3559;
  assign T_166_up_idx = T_3527;
  assign T_166_up_done = T_3528;
  assign T_166_down_idx = 3'h0;
  assign T_166_down_done = T_3529;
  assign T_186_pending = T_3161;
  assign T_186_up_idx = T_3102;
  assign T_186_up_done = T_3103;
  assign T_186_down_idx = T_3144;
  assign T_186_down_done = T_3145;
  assign T_210_pending = T_2976;
  assign T_210_up_idx = T_2919;
  assign T_210_up_done = T_2920;
  assign T_210_down_idx = T_2959;
  assign T_210_down_done = T_2960;
  assign GEN_432 = {{7'd0}, 1'h0};
  assign T_219 = T_201 != GEN_432;
  assign T_220 = T_199 | T_219;
  assign T_221 = T_220 | T_210_pending;
  assign T_247_sharers = 1'h0;
  assign T_299_state = {{1'd0}, 1'h0};
  assign T_395_inner_sharers = T_247_sharers;
  assign T_395_outer_state = T_299_state;
  assign T_1733 = T_55 == 4'h0;
  assign T_1734 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1735 = T_1733 & T_1734;
  assign T_1736 = T_1735 & io_alloc_iacq_should;
  assign T_1745_0 = 3'h3;
  assign T_1747 = T_1745_0 == io_inner_acquire_bits_a_type;
  assign T_1750 = io_inner_acquire_bits_is_builtin_type & T_1747;
  assign T_1751 = T_1736 & T_1750;
  assign T_1760_0 = 3'h3;
  assign T_1762 = T_1760_0 == io_inner_acquire_bits_a_type;
  assign T_1765 = io_inner_acquire_bits_is_builtin_type & T_1762;
  assign T_1767 = T_1765 == 1'h0;
  assign GEN_433 = {{2'd0}, 1'h0};
  assign T_1769 = io_inner_acquire_bits_addr_beat == GEN_433;
  assign T_1770 = T_1767 | T_1769;
  assign T_1772 = T_1770 == 1'h0;
  assign T_1773 = T_1751 & T_1772;
  assign T_1775 = T_1773 == 1'h0;
  assign T_1776 = T_1775 | reset;
  assign T_1778 = T_1776 == 1'h0;
  assign T_1779 = T_55 != 4'h0;
  assign T_1780 = T_1779 & T_153;
  assign T_1782 = T_99_a_type == 3'h5;
  assign T_1784 = T_99_a_type == 3'h6;
  assign T_1785 = T_1782 | T_1784;
  assign T_1786 = T_99_is_builtin_type & T_1785;
  assign T_1787 = T_1780 & T_1786;
  assign T_1789 = T_1787 == 1'h0;
  assign T_1790 = T_1789 | reset;
  assign T_1792 = T_1790 == 1'h0;
  assign T_1796 = T_99_a_type == 3'h4;
  assign T_1797 = T_99_is_builtin_type & T_1796;
  assign T_1798 = T_1780 & T_1797;
  assign T_1800 = T_1798 == 1'h0;
  assign T_1801 = T_1800 | reset;
  assign T_1803 = T_1801 == 1'h0;
  assign T_1817_0 = 64'h0;
  assign T_1817_1 = 64'h0;
  assign T_1817_2 = 64'h0;
  assign T_1817_3 = 64'h0;
  assign T_1817_4 = 64'h0;
  assign T_1817_5 = 64'h0;
  assign T_1817_6 = 64'h0;
  assign T_1817_7 = 64'h0;
  assign T_1835_0 = 8'h0;
  assign T_1835_1 = 8'h0;
  assign T_1835_2 = 8'h0;
  assign T_1835_3 = 8'h0;
  assign T_1835_4 = 8'h0;
  assign T_1835_5 = 8'h0;
  assign T_1835_6 = 8'h0;
  assign T_1835_7 = 8'h0;
  assign T_1841 = io_inner_acquire_bits_addr_block == T_57;
  assign T_1842 = T_1779 & T_1841;
  assign T_1844 = io_inner_release_bits_addr_block == T_57;
  assign T_1845 = T_1779 & T_1844;
  assign T_1847 = io_outer_probe_bits_addr_block == T_57;
  assign T_1848 = T_1779 & T_1847;
  assign Queue_14_1_clk = clk;
  assign Queue_14_1_reset = reset;
  assign Queue_14_1_io_enq_valid = T_1929;
  assign Queue_14_1_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign Queue_14_1_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign Queue_14_1_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign Queue_14_1_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign Queue_14_1_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign Queue_14_1_io_deq_ready = GEN_349;
  assign T_1884 = T_1733 & io_alloc_iacq_should;
  assign T_1885 = T_1884 & io_inner_acquire_valid;
  assign T_1887 = T_99_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1896_0 = 3'h3;
  assign T_1898 = T_1896_0 == T_99_a_type;
  assign T_1901 = T_99_is_builtin_type & T_1898;
  assign T_1902 = T_1887 & T_1901;
  assign T_1903 = T_1902 & T_153;
  assign T_1904 = T_175 >> io_inner_acquire_bits_addr_beat;
  assign T_1905 = T_1904[0];
  assign T_1906 = T_1903 & T_1905;
  assign T_1908 = T_1906 & io_inner_acquire_valid;
  assign T_1917_0 = 3'h3;
  assign T_1919 = T_1917_0 == io_inner_acquire_bits_a_type;
  assign T_1922 = io_inner_acquire_bits_is_builtin_type & T_1919;
  assign T_1924 = T_1922 == 1'h0;
  assign T_1927 = T_1924 | T_1769;
  assign T_1928 = T_1908 & T_1927;
  assign T_1929 = T_1885 | T_1928;
  assign T_1930_client_xact_id = Queue_14_1_io_deq_valid ? Queue_14_1_io_deq_bits_client_xact_id : Queue_14_1_io_enq_bits_client_xact_id;
  assign T_1930_addr_beat = Queue_14_1_io_deq_valid ? Queue_14_1_io_deq_bits_addr_beat : Queue_14_1_io_enq_bits_addr_beat;
  assign T_1930_client_id = Queue_14_1_io_deq_valid ? Queue_14_1_io_deq_bits_client_id : Queue_14_1_io_enq_bits_client_id;
  assign T_1930_is_builtin_type = Queue_14_1_io_deq_valid ? Queue_14_1_io_deq_bits_is_builtin_type : Queue_14_1_io_enq_bits_is_builtin_type;
  assign T_1930_a_type = Queue_14_1_io_deq_valid ? Queue_14_1_io_deq_bits_a_type : Queue_14_1_io_enq_bits_a_type;
  assign GEN_435 = {{1'd0}, 1'h0};
  assign T_1960 = Queue_14_1_io_count > GEN_435;
  assign T_1962 = T_1779 | io_alloc_iacq_should;
  assign T_1972_0 = 3'h2;
  assign T_1972_1 = 3'h3;
  assign T_1972_2 = 3'h4;
  assign T_1974 = T_1972_0 == io_inner_acquire_bits_a_type;
  assign T_1975 = T_1972_1 == io_inner_acquire_bits_a_type;
  assign T_1976 = T_1972_2 == io_inner_acquire_bits_a_type;
  assign T_1979 = T_1974 | T_1975;
  assign T_1980 = T_1979 | T_1976;
  assign T_1981 = io_inner_acquire_bits_is_builtin_type & T_1980;
  assign T_1982 = T_1734 & T_1981;
  assign GEN_436 = {{7'd0}, T_1982};
  assign T_1984 = 8'h0 - GEN_436;
  assign T_1985 = T_1984[7:0];
  assign T_1986 = ~ T_1985;
  assign GEN_437 = {{7'd0}, 1'h1};
  assign T_1988 = GEN_437 << io_inner_acquire_bits_addr_beat;
  assign T_1989 = ~ T_1988;
  assign T_1990 = T_1986 | T_1989;
  assign T_1991 = T_175 & T_1990;
  assign T_2001_0 = 3'h3;
  assign T_2003 = T_2001_0 == io_inner_acquire_bits_a_type;
  assign T_2006 = io_inner_acquire_bits_is_builtin_type & T_2003;
  assign T_2007 = T_1734 & T_2006;
  assign T_2010 = T_2007 & T_1769;
  assign T_2019 = T_2010 ? 8'hfe : 8'h0;
  assign T_2020 = T_1991 | T_2019;
  assign GEN_32 = T_1962 ? T_2020 : T_175;
  assign GEN_439 = {{3'd0}, 1'h0};
  assign T_2028 = 4'h8 * GEN_439;
  assign T_2030 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_2031 = io_inner_acquire_bits_is_builtin_type & T_2030;
  assign T_2033 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_2034 = io_inner_acquire_bits_is_builtin_type & T_2033;
  assign T_2035 = T_2031 | T_2034;
  assign T_2036 = io_inner_acquire_bits_union[5:1];
  assign T_2037 = T_2035 ? 5'h1 : T_2036;
  assign T_2038 = io_inner_acquire_bits_union[11:9];
  assign T_2039 = io_inner_acquire_bits_union[8:6];
  assign T_2052_0 = 3'h2;
  assign T_2052_1 = 3'h3;
  assign T_2052_2 = 3'h4;
  assign T_2054 = T_2052_0 == io_inner_acquire_bits_a_type;
  assign T_2055 = T_2052_1 == io_inner_acquire_bits_a_type;
  assign T_2056 = T_2052_2 == io_inner_acquire_bits_a_type;
  assign T_2059 = T_2054 | T_2055;
  assign T_2060 = T_2059 | T_2056;
  assign T_2061 = io_inner_acquire_bits_is_builtin_type & T_2060;
  assign T_2062 = T_1734 & T_2061;
  assign GEN_440 = {{7'd0}, T_2062};
  assign T_2064 = 8'h0 - GEN_440;
  assign T_2065 = T_2064[7:0];
  assign T_2066 = ~ T_2065;
  assign T_2070 = T_2066 | T_1989;
  assign T_2072 = T_2034 ? T_2070 : {{7'd0}, 1'h0};
  assign GEN_33 = T_1885 ? io_inner_acquire_bits_addr_block : T_57;
  assign GEN_34 = T_1885 ? 1'h0 : T_59;
  assign GEN_35 = T_1885 ? T_2028 : T_61;
  assign GEN_36 = T_1885 ? T_2037 : T_63;
  assign GEN_37 = T_1885 ? T_2038 : T_65;
  assign GEN_38 = T_1885 ? T_2039 : T_67;
  assign GEN_42 = T_1885 ? T_2072 : GEN_32;
  assign GEN_43 = T_1885 ? {{7'd0}, 1'h0} : T_177;
  assign GEN_44 = T_1885 ? 4'h5 : T_55;
  assign T_2075 = T_175 != GEN_432;
  assign T_2088_0 = 3'h3;
  assign T_2090 = T_2088_0 == T_99_a_type;
  assign T_2093 = T_99_is_builtin_type & T_2090;
  assign T_2094 = T_1887 & T_2093;
  assign T_2095 = T_2094 & T_153;
  assign T_2098 = T_2095 & T_1905;
  assign T_2099 = T_1733 | T_2098;
  assign T_2100 = ~ T_177;
  assign skip_outer_acquire = T_2100 == GEN_432;
  assign T_2109 = 3'h4 == T_99_a_type;
  assign T_2110 = T_2109 ? 2'h0 : 2'h2;
  assign T_2111 = 3'h6 == T_99_a_type;
  assign T_2112 = T_2111 ? 2'h0 : T_2110;
  assign T_2113 = 3'h5 == T_99_a_type;
  assign T_2114 = T_2113 ? 2'h2 : T_2112;
  assign T_2115 = 3'h2 == T_99_a_type;
  assign T_2116 = T_2115 ? 2'h0 : T_2114;
  assign T_2117 = 3'h0 == T_99_a_type;
  assign T_2118 = T_2117 ? 2'h2 : T_2116;
  assign T_2119 = 3'h3 == T_99_a_type;
  assign T_2120 = T_2119 ? 2'h0 : T_2118;
  assign T_2121 = 3'h1 == T_99_a_type;
  assign T_2122 = T_2121 ? 2'h2 : T_2120;
  assign GEN_444 = {{2'd0}, 1'h1};
  assign T_2123 = GEN_444 == T_99_a_type;
  assign T_2124 = T_2123 ? 2'h0 : 2'h2;
  assign T_2125 = GEN_433 == T_99_a_type;
  assign T_2126 = T_2125 ? 2'h1 : T_2124;
  assign T_2127 = T_99_is_builtin_type ? T_2122 : T_2126;
  assign T_2155_addr_block = T_57;
  assign T_2155_p_type = T_2127;
  assign T_2155_client_id = 1'h0;
  assign T_2183 = skip_outer_acquire == 1'h0;
  assign T_2184 = T_2183 ? 4'h6 : 4'h7;
  assign T_2193_pending = T_2276;
  assign T_2193_up_idx = 3'h0;
  assign T_2193_up_done = T_2201;
  assign T_2193_down_idx = T_2259;
  assign T_2193_down_done = T_2260;
  assign T_2201 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2202 = ~ T_2201;
  assign GEN_446 = {{1'd0}, 1'h1};
  assign T_2204 = GEN_446 << io_inner_probe_bits_client_id;
  assign T_2205 = ~ T_2204;
  assign GEN_447 = {{1'd0}, T_2202};
  assign T_2206 = GEN_447 | T_2205;
  assign GEN_448 = {{1'd0}, T_195};
  assign T_2207 = GEN_448 & T_2206;
  assign T_2208 = T_55 == 4'h5;
  assign T_2211 = T_2208 & T_195;
  assign T_2228 = io_inner_release_ready & io_inner_release_valid;
  assign T_2231 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2232 = T_1779 & T_2231;
  assign T_2233 = T_2228 & T_2232;
  assign T_2240_0 = 3'h0;
  assign T_2240_1 = 3'h1;
  assign T_2240_2 = 3'h2;
  assign T_2242 = T_2240_0 == io_inner_release_bits_r_type;
  assign T_2243 = T_2240_1 == io_inner_release_bits_r_type;
  assign T_2244 = T_2240_2 == io_inner_release_bits_r_type;
  assign T_2247 = T_2242 | T_2243;
  assign T_2248 = T_2247 | T_2244;
  assign T_2250 = T_2233 & T_2248;
  assign T_2254 = T_2252 == 3'h7;
  assign T_2256 = T_2252 + GEN_444;
  assign T_2257 = T_2256[2:0];
  assign GEN_46 = T_2250 ? T_2257 : T_2252;
  assign T_2258 = T_2250 & T_2254;
  assign T_2259 = T_2248 ? T_2252 : {{2'd0}, 1'h0};
  assign T_2260 = T_2248 ? T_2258 : T_2233;
  assign T_2264 = T_2260 == 1'h0;
  assign T_2265 = T_2201 & T_2264;
  assign T_2267 = T_2262 + 1'h1;
  assign T_2268 = T_2267[0:0];
  assign GEN_47 = T_2265 ? T_2268 : T_2262;
  assign T_2270 = T_2201 == 1'h0;
  assign T_2271 = T_2260 & T_2270;
  assign T_2273 = T_2262 - 1'h1;
  assign T_2274 = T_2273[0:0];
  assign GEN_48 = T_2271 ? T_2274 : GEN_47;
  assign T_2276 = T_2262 > 1'h0;
  assign T_2280 = T_195 | T_2193_pending;
  assign T_2282 = T_2280 == 1'h0;
  assign T_2283 = T_2208 & T_2282;
  assign GEN_49 = T_2283 ? T_2184 : GEN_44;
  assign T_2287 = T_1733 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2288 = T_2287 & io_inner_release_bits_voluntary;
  assign T_2293 = T_2228 & T_2288;
  assign T_2300_0 = 3'h0;
  assign T_2300_1 = 3'h1;
  assign T_2300_2 = 3'h2;
  assign T_2302 = T_2300_0 == io_inner_release_bits_r_type;
  assign T_2303 = T_2300_1 == io_inner_release_bits_r_type;
  assign T_2304 = T_2300_2 == io_inner_release_bits_r_type;
  assign T_2307 = T_2302 | T_2303;
  assign T_2308 = T_2307 | T_2304;
  assign T_2310 = T_2293 & T_2308;
  assign T_2314 = T_2312 == 3'h7;
  assign T_2316 = T_2312 + GEN_444;
  assign T_2317 = T_2316[2:0];
  assign GEN_50 = T_2310 ? T_2317 : T_2312;
  assign T_2318 = T_2310 & T_2314;
  assign T_2319 = T_2308 ? T_2312 : {{2'd0}, 1'h0};
  assign T_2320 = T_2308 ? T_2318 : T_2293;
  assign T_2321 = io_inner_grant_ready & io_inner_grant_valid;
  assign GEN_452 = {{1'd0}, 3'h0};
  assign T_2324 = io_inner_grant_bits_g_type == GEN_452;
  assign T_2325 = io_inner_grant_bits_is_builtin_type & T_2324;
  assign T_2326 = T_1779 & T_2325;
  assign T_2327 = T_2321 & T_2326;
  assign T_2335_0 = 3'h5;
  assign GEN_453 = {{1'd0}, T_2335_0};
  assign T_2337 = GEN_453 == io_inner_grant_bits_g_type;
  assign T_2345_0 = 2'h0;
  assign T_2345_1 = 2'h1;
  assign GEN_454 = {{2'd0}, T_2345_0};
  assign T_2347 = GEN_454 == io_inner_grant_bits_g_type;
  assign GEN_455 = {{2'd0}, T_2345_1};
  assign T_2348 = GEN_455 == io_inner_grant_bits_g_type;
  assign T_2351 = T_2347 | T_2348;
  assign T_2352 = io_inner_grant_bits_is_builtin_type ? T_2337 : T_2351;
  assign T_2354 = T_2327 & T_2352;
  assign T_2358 = T_2356 == 3'h7;
  assign T_2360 = T_2356 + GEN_444;
  assign T_2361 = T_2360[2:0];
  assign GEN_51 = T_2354 ? T_2361 : T_2356;
  assign T_2362 = T_2354 & T_2358;
  assign T_2363 = T_2352 ? T_2356 : {{2'd0}, 1'h0};
  assign T_2364 = T_2352 ? T_2362 : T_2327;
  assign T_2368 = T_2364 == 1'h0;
  assign T_2369 = T_2320 & T_2368;
  assign T_2371 = T_2366 + 1'h1;
  assign T_2372 = T_2371[0:0];
  assign GEN_52 = T_2369 ? T_2372 : T_2366;
  assign T_2374 = T_2320 == 1'h0;
  assign T_2375 = T_2364 & T_2374;
  assign T_2377 = T_2366 - 1'h1;
  assign T_2378 = T_2377[0:0];
  assign GEN_53 = T_2375 ? T_2378 : GEN_52;
  assign T_2380 = T_2366 > 1'h0;
  assign T_2382 = T_1733 & io_alloc_irel_should;
  assign T_2383 = T_2382 & io_inner_release_valid;
  assign GEN_54 = T_2383 ? io_inner_release_bits_addr_block : GEN_33;
  assign GEN_55 = T_2383 ? 4'h7 : GEN_49;
  assign T_2386 = T_1844 & io_inner_release_bits_voluntary;
  assign T_2392_0 = 4'h0;
  assign T_2392_1 = 4'h8;
  assign T_2394 = T_2392_0 == T_55;
  assign T_2395 = T_2392_1 == T_55;
  assign T_2398 = T_2394 | T_2395;
  assign T_2400 = T_2398 == 1'h0;
  assign T_2401 = T_2386 & T_2400;
  assign T_2403 = T_44 == 1'h0;
  assign T_2404 = T_2401 & T_2403;
  assign T_2405 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2407 = T_2405 == 1'h0;
  assign T_2408 = T_2404 & T_2407;
  assign T_2411 = T_2321 == 1'h0;
  assign T_2412 = T_2408 & T_2411;
  assign T_2414 = T_144_pending == 1'h0;
  assign T_2415 = T_2412 & T_2414;
  assign T_2422_0 = 3'h0;
  assign T_2422_1 = 3'h1;
  assign T_2422_2 = 3'h2;
  assign T_2424 = T_2422_0 == io_inner_release_bits_r_type;
  assign T_2425 = T_2422_1 == io_inner_release_bits_r_type;
  assign T_2426 = T_2422_2 == io_inner_release_bits_r_type;
  assign T_2429 = T_2424 | T_2425;
  assign T_2430 = T_2429 | T_2426;
  assign T_2433 = T_2430 == 1'h0;
  assign T_2435 = io_inner_release_bits_addr_beat == GEN_433;
  assign T_2436 = T_2433 | T_2435;
  assign T_2437 = T_2415 & T_2436;
  assign T_2438 = io_alloc_irel_should | T_2437;
  assign T_2445_0 = 3'h0;
  assign T_2445_1 = 3'h1;
  assign T_2445_2 = 3'h2;
  assign T_2447 = T_2445_0 == io_inner_release_bits_r_type;
  assign T_2448 = T_2445_1 == io_inner_release_bits_r_type;
  assign T_2449 = T_2445_2 == io_inner_release_bits_r_type;
  assign T_2452 = T_2447 | T_2448;
  assign T_2453 = T_2452 | T_2449;
  assign T_2461_0 = 3'h0;
  assign T_2461_1 = 3'h1;
  assign T_2461_2 = 3'h2;
  assign T_2463 = T_2461_0 == io_inner_release_bits_r_type;
  assign T_2464 = T_2461_1 == io_inner_release_bits_r_type;
  assign T_2465 = T_2461_2 == io_inner_release_bits_r_type;
  assign T_2468 = T_2463 | T_2464;
  assign T_2469 = T_2468 | T_2465;
  assign T_2470 = T_2228 & T_2469;
  assign GEN_458 = {{7'd0}, T_2470};
  assign T_2472 = 8'h0 - GEN_458;
  assign T_2473 = T_2472[7:0];
  assign T_2474 = ~ T_2473;
  assign T_2476 = GEN_437 << io_inner_release_bits_addr_beat;
  assign T_2477 = ~ T_2476;
  assign T_2478 = T_2474 | T_2477;
  assign T_2480 = T_2453 ? T_2478 : {{7'd0}, 1'h0};
  assign GEN_56 = T_2438 ? io_inner_release_bits_r_type : T_129;
  assign GEN_57 = T_2438 ? io_inner_release_bits_client_id : T_131;
  assign GEN_58 = T_2438 ? io_inner_release_bits_client_xact_id : T_133;
  assign GEN_65 = T_2438 ? T_2480 : T_135;
  assign T_2484 = T_1844 & T_2231;
  assign T_2486 = T_2484 & T_2208;
  assign T_2488 = T_2438 == 1'h0;
  assign T_2489 = T_2488 & T_2486;
  assign T_2496_0 = 3'h0;
  assign T_2496_1 = 3'h1;
  assign T_2496_2 = 3'h2;
  assign T_2498 = T_2496_0 == io_inner_release_bits_r_type;
  assign T_2499 = T_2496_1 == io_inner_release_bits_r_type;
  assign T_2500 = T_2496_2 == io_inner_release_bits_r_type;
  assign T_2503 = T_2498 | T_2499;
  assign T_2504 = T_2503 | T_2500;
  assign T_2505 = T_2228 & T_2504;
  assign GEN_460 = {{7'd0}, T_2505};
  assign T_2507 = 8'h0 - GEN_460;
  assign T_2508 = T_2507[7:0];
  assign T_2509 = ~ T_2508;
  assign T_2513 = T_2509 | T_2477;
  assign T_2514 = T_135 & T_2513;
  assign GEN_69 = T_2489 ? T_2514 : GEN_65;
  assign GEN_75 = T_2228 ? GEN_56 : T_129;
  assign GEN_76 = T_2228 ? GEN_57 : T_131;
  assign GEN_77 = T_2228 ? GEN_58 : T_133;
  assign GEN_84 = T_2228 ? GEN_69 : T_135;
  assign T_2520_0 = 4'h3;
  assign T_2520_1 = 4'h4;
  assign T_2520_2 = 4'h5;
  assign T_2520_3 = 4'h7;
  assign T_2522 = T_2520_0 == T_55;
  assign T_2523 = T_2520_1 == T_55;
  assign T_2524 = T_2520_2 == T_55;
  assign T_2525 = T_2520_3 == T_55;
  assign T_2528 = T_2522 | T_2523;
  assign T_2529 = T_2528 | T_2524;
  assign T_2530 = T_2529 | T_2525;
  assign T_2531 = T_2530 & T_144_pending;
  assign T_2533 = T_135 != GEN_432;
  assign T_2534 = T_2533 | T_210_pending;
  assign T_2536 = T_2534 == 1'h0;
  assign T_2537 = T_2531 & T_2536;
  assign T_2572_addr_beat = {{2'd0}, 1'h0};
  assign T_2572_addr_block = T_57;
  assign T_2572_client_xact_id = T_133;
  assign T_2572_voluntary = 1'h1;
  assign T_2572_r_type = T_129;
  assign T_2572_data = {{63'd0}, 1'h0};
  assign T_2572_client_id = T_131;
  assign T_2639_addr_beat = {{2'd0}, 1'h0};
  assign T_2639_client_xact_id = T_2572_client_xact_id;
  assign T_2639_manager_xact_id = {{2'd0}, 1'h0};
  assign T_2639_is_builtin_type = 1'h1;
  assign T_2639_g_type = {{1'd0}, 3'h0};
  assign T_2639_data = {{63'd0}, 1'h0};
  assign T_2639_client_id = T_2572_client_id;
  assign T_2679_0 = 4'h0;
  assign T_2679_1 = 4'h8;
  assign T_2681 = T_2679_0 == T_55;
  assign T_2682 = T_2679_1 == T_55;
  assign T_2685 = T_2681 | T_2682;
  assign T_2687 = T_2685 == 1'h0;
  assign T_2688 = T_2386 & T_2687;
  assign T_2691 = T_2688 & T_2403;
  assign T_2695 = T_2691 & T_2407;
  assign T_2699 = T_2695 & T_2411;
  assign T_2702 = T_2699 & T_2414;
  assign T_2709 = T_2702 | T_2486;
  assign T_2716_0 = 3'h0;
  assign T_2716_1 = 3'h1;
  assign T_2716_2 = 3'h2;
  assign T_2718 = T_2716_0 == io_inner_release_bits_r_type;
  assign T_2719 = T_2716_1 == io_inner_release_bits_r_type;
  assign T_2720 = T_2716_2 == io_inner_release_bits_r_type;
  assign T_2723 = T_2718 | T_2719;
  assign T_2724 = T_2723 | T_2720;
  assign T_2725 = T_2228 & T_2724;
  assign GEN_0 = GEN_94;
  assign GEN_88 = GEN_444 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_465 = {{1'd0}, 2'h2};
  assign GEN_89 = GEN_465 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_88;
  assign GEN_466 = {{1'd0}, 2'h3};
  assign GEN_90 = GEN_466 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_89;
  assign GEN_91 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_90;
  assign GEN_92 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_91;
  assign GEN_93 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_92;
  assign GEN_94 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_93;
  assign T_2726 = GEN_0[0];
  assign GEN_1 = GEN_94;
  assign T_2727 = GEN_1[1];
  assign GEN_2 = GEN_94;
  assign T_2728 = GEN_2[2];
  assign GEN_3 = GEN_94;
  assign T_2729 = GEN_3[3];
  assign GEN_4 = GEN_94;
  assign T_2730 = GEN_4[4];
  assign GEN_5 = GEN_94;
  assign T_2731 = GEN_5[5];
  assign GEN_6 = GEN_94;
  assign T_2732 = GEN_6[6];
  assign GEN_7 = GEN_94;
  assign T_2733 = GEN_7[7];
  assign GEN_488 = {{7'd0}, T_2726};
  assign T_2735 = 8'h0 - GEN_488;
  assign T_2736 = T_2735[7:0];
  assign GEN_489 = {{7'd0}, T_2727};
  assign T_2738 = 8'h0 - GEN_489;
  assign T_2739 = T_2738[7:0];
  assign GEN_490 = {{7'd0}, T_2728};
  assign T_2741 = 8'h0 - GEN_490;
  assign T_2742 = T_2741[7:0];
  assign GEN_491 = {{7'd0}, T_2729};
  assign T_2744 = 8'h0 - GEN_491;
  assign T_2745 = T_2744[7:0];
  assign GEN_492 = {{7'd0}, T_2730};
  assign T_2747 = 8'h0 - GEN_492;
  assign T_2748 = T_2747[7:0];
  assign GEN_493 = {{7'd0}, T_2731};
  assign T_2750 = 8'h0 - GEN_493;
  assign T_2751 = T_2750[7:0];
  assign GEN_494 = {{7'd0}, T_2732};
  assign T_2753 = 8'h0 - GEN_494;
  assign T_2754 = T_2753[7:0];
  assign GEN_495 = {{7'd0}, T_2733};
  assign T_2756 = 8'h0 - GEN_495;
  assign T_2757 = T_2756[7:0];
  assign T_2763_0 = T_2736;
  assign T_2763_1 = T_2739;
  assign T_2763_2 = T_2742;
  assign T_2763_3 = T_2745;
  assign T_2763_4 = T_2748;
  assign T_2763_5 = T_2751;
  assign T_2763_6 = T_2754;
  assign T_2763_7 = T_2757;
  assign T_2765 = {T_2763_1,T_2763_0};
  assign T_2766 = {T_2763_3,T_2763_2};
  assign T_2767 = {T_2766,T_2765};
  assign T_2768 = {T_2763_5,T_2763_4};
  assign T_2769 = {T_2763_7,T_2763_6};
  assign T_2770 = {T_2769,T_2768};
  assign T_2771 = {T_2770,T_2767};
  assign T_2772 = ~ T_2771;
  assign T_2773 = T_2772 & io_inner_release_bits_data;
  assign GEN_8 = GEN_150;
  assign GEN_144 = GEN_444 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_145 = GEN_465 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_144;
  assign GEN_146 = GEN_466 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_145;
  assign GEN_147 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_146;
  assign GEN_148 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_147;
  assign GEN_149 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_148;
  assign GEN_150 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_149;
  assign T_2774 = T_2771 & GEN_8;
  assign T_2775 = T_2773 | T_2774;
  assign GEN_9 = T_2775;
  assign GEN_151 = GEN_433 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_152 = GEN_444 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_153 = GEN_465 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_154 = GEN_466 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_155 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_156 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_157 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_158 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_177 = T_2725 ? GEN_151 : data_buffer_0;
  assign GEN_178 = T_2725 ? GEN_152 : data_buffer_1;
  assign GEN_179 = T_2725 ? GEN_153 : data_buffer_2;
  assign GEN_180 = T_2725 ? GEN_154 : data_buffer_3;
  assign GEN_181 = T_2725 ? GEN_155 : data_buffer_4;
  assign GEN_182 = T_2725 ? GEN_156 : data_buffer_5;
  assign GEN_183 = T_2725 ? GEN_157 : data_buffer_6;
  assign GEN_184 = T_2725 ? GEN_158 : data_buffer_7;
  assign T_2806_state = 2'h2;
  assign T_2832 = T_1779 | io_alloc_irel_should;
  assign T_2833 = io_outer_release_ready & io_outer_release_valid;
  assign T_2839_0 = 3'h0;
  assign T_2839_1 = 3'h1;
  assign T_2839_2 = 3'h2;
  assign T_2841 = T_2839_0 == io_outer_release_bits_r_type;
  assign T_2842 = T_2839_1 == io_outer_release_bits_r_type;
  assign T_2843 = T_2839_2 == io_outer_release_bits_r_type;
  assign T_2846 = T_2841 | T_2842;
  assign T_2847 = T_2846 | T_2843;
  assign T_2848 = T_2833 & T_2847;
  assign GEN_503 = {{7'd0}, T_2848};
  assign T_2850 = 8'h0 - GEN_503;
  assign T_2851 = T_2850[7:0];
  assign T_2852 = ~ T_2851;
  assign T_2854 = GEN_437 << io_outer_release_bits_addr_beat;
  assign T_2855 = ~ T_2854;
  assign T_2856 = T_2852 | T_2855;
  assign T_2857 = T_201 & T_2856;
  assign T_2865_0 = 3'h0;
  assign T_2865_1 = 3'h1;
  assign T_2865_2 = 3'h2;
  assign T_2867 = T_2865_0 == io_inner_release_bits_r_type;
  assign T_2868 = T_2865_1 == io_inner_release_bits_r_type;
  assign T_2869 = T_2865_2 == io_inner_release_bits_r_type;
  assign T_2872 = T_2867 | T_2868;
  assign T_2873 = T_2872 | T_2869;
  assign T_2874 = T_2228 & T_2873;
  assign GEN_505 = {{7'd0}, T_2874};
  assign T_2877 = 8'h0 - GEN_505;
  assign T_2878 = T_2877[7:0];
  assign T_2881 = T_2878 & T_2476;
  assign T_2882 = T_2857 | T_2881;
  assign T_2883 = T_2882 | GEN_432;
  assign GEN_191 = T_2832 ? T_2883 : T_201;
  assign GEN_193 = T_2833 ? 1'h0 : T_199;
  assign T_2893 = T_2833 & io_outer_release_bits_voluntary;
  assign T_2900_0 = 3'h0;
  assign T_2900_1 = 3'h1;
  assign T_2900_2 = 3'h2;
  assign T_2902 = T_2900_0 == io_outer_release_bits_r_type;
  assign T_2903 = T_2900_1 == io_outer_release_bits_r_type;
  assign T_2904 = T_2900_2 == io_outer_release_bits_r_type;
  assign T_2907 = T_2902 | T_2903;
  assign T_2908 = T_2907 | T_2904;
  assign T_2910 = T_2893 & T_2908;
  assign T_2914 = T_2912 == 3'h7;
  assign T_2916 = T_2912 + GEN_444;
  assign T_2917 = T_2916[2:0];
  assign GEN_194 = T_2910 ? T_2917 : T_2912;
  assign T_2918 = T_2910 & T_2914;
  assign T_2919 = T_2908 ? T_2912 : {{2'd0}, 1'h0};
  assign T_2920 = T_2908 ? T_2918 : T_2893;
  assign T_2923 = io_outer_grant_bits_g_type == GEN_452;
  assign T_2924 = io_outer_grant_bits_is_builtin_type & T_2923;
  assign T_2925 = T_2405 & T_2924;
  assign T_2933_0 = 3'h5;
  assign GEN_510 = {{1'd0}, T_2933_0};
  assign T_2935 = GEN_510 == io_outer_grant_bits_g_type;
  assign T_2943_0 = 1'h0;
  assign GEN_511 = {{3'd0}, T_2943_0};
  assign T_2945 = GEN_511 == io_outer_grant_bits_g_type;
  assign T_2948 = io_outer_grant_bits_is_builtin_type ? T_2935 : T_2945;
  assign T_2950 = T_2925 & T_2948;
  assign T_2954 = T_2952 == 3'h7;
  assign T_2956 = T_2952 + GEN_444;
  assign T_2957 = T_2956[2:0];
  assign GEN_195 = T_2950 ? T_2957 : T_2952;
  assign T_2958 = T_2950 & T_2954;
  assign T_2959 = T_2948 ? T_2952 : {{2'd0}, 1'h0};
  assign T_2960 = T_2948 ? T_2958 : T_2925;
  assign T_2964 = T_2960 == 1'h0;
  assign T_2965 = T_2920 & T_2964;
  assign T_2967 = T_2962 + 1'h1;
  assign T_2968 = T_2967[0:0];
  assign GEN_196 = T_2965 ? T_2968 : T_2962;
  assign T_2970 = T_2920 == 1'h0;
  assign T_2971 = T_2960 & T_2970;
  assign T_2973 = T_2962 - 1'h1;
  assign T_2974 = T_2973[0:0];
  assign GEN_197 = T_2971 ? T_2974 : GEN_196;
  assign T_2976 = T_2962 > 1'h0;
  assign T_2977 = T_55 == 4'h7;
  assign T_2983_0 = 3'h0;
  assign T_2983_1 = 3'h1;
  assign T_2983_2 = 3'h2;
  assign T_2985 = T_2983_0 == io_outer_release_bits_r_type;
  assign T_2986 = T_2983_1 == io_outer_release_bits_r_type;
  assign T_2987 = T_2983_2 == io_outer_release_bits_r_type;
  assign T_2990 = T_2985 | T_2986;
  assign T_2991 = T_2990 | T_2987;
  assign T_2992 = T_201 >> T_210_up_idx;
  assign T_2993 = T_2992[0];
  assign T_2995 = T_2991 ? T_2993 : T_221;
  assign T_2996 = T_2977 & T_2995;
  assign T_3004_0 = 2'h2;
  assign T_3006 = T_3004_0 == T_2806_state;
  assign T_3009 = T_3006 ? 3'h0 : 3'h3;
  assign T_3045_addr_beat = T_210_up_idx;
  assign T_3045_addr_block = T_57;
  assign T_3045_client_xact_id = {{2'd0}, 1'h0};
  assign T_3045_voluntary = 1'h1;
  assign T_3045_r_type = T_3009;
  assign T_3045_data = GEN_10;
  assign GEN_10 = GEN_204;
  assign GEN_198 = GEN_444 == T_210_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_199 = GEN_465 == T_210_up_idx ? data_buffer_2 : GEN_198;
  assign GEN_200 = GEN_466 == T_210_up_idx ? data_buffer_3 : GEN_199;
  assign GEN_201 = 3'h4 == T_210_up_idx ? data_buffer_4 : GEN_200;
  assign GEN_202 = 3'h5 == T_210_up_idx ? data_buffer_5 : GEN_201;
  assign GEN_203 = 3'h6 == T_210_up_idx ? data_buffer_6 : GEN_202;
  assign GEN_204 = 3'h7 == T_210_up_idx ? data_buffer_7 : GEN_203;
  assign T_3074 = T_99_is_builtin_type == 1'h0;
  assign T_3076 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_3087_0 = 3'h3;
  assign T_3089 = T_3087_0 == io_outer_acquire_bits_a_type;
  assign T_3092 = io_outer_acquire_bits_is_builtin_type & T_3089;
  assign T_3093 = T_3076 & T_3092;
  assign T_3097 = T_3095 == 3'h7;
  assign T_3099 = T_3095 + GEN_444;
  assign T_3100 = T_3099[2:0];
  assign GEN_205 = T_3093 ? T_3100 : T_3095;
  assign T_3101 = T_3093 & T_3097;
  assign T_3102 = T_3092 ? T_3095 : T_69;
  assign T_3103 = T_3092 ? T_3101 : T_3076;
  assign T_3109 = T_2924 == 1'h0;
  assign T_3110 = T_2405 & T_3109;
  assign T_3118_0 = 3'h5;
  assign GEN_518 = {{1'd0}, T_3118_0};
  assign T_3120 = GEN_518 == io_outer_grant_bits_g_type;
  assign T_3128_0 = 1'h0;
  assign GEN_519 = {{3'd0}, T_3128_0};
  assign T_3130 = GEN_519 == io_outer_grant_bits_g_type;
  assign T_3133 = io_outer_grant_bits_is_builtin_type ? T_3120 : T_3130;
  assign T_3135 = T_3110 & T_3133;
  assign T_3139 = T_3137 == 3'h7;
  assign T_3141 = T_3137 + GEN_444;
  assign T_3142 = T_3141[2:0];
  assign GEN_206 = T_3135 ? T_3142 : T_3137;
  assign T_3143 = T_3135 & T_3139;
  assign T_3144 = T_3133 ? T_3137 : T_69;
  assign T_3145 = T_3133 ? T_3143 : T_3110;
  assign T_3149 = T_3145 == 1'h0;
  assign T_3150 = T_3103 & T_3149;
  assign T_3152 = T_3147 + 1'h1;
  assign T_3153 = T_3152[0:0];
  assign GEN_207 = T_3150 ? T_3153 : T_3147;
  assign T_3155 = T_3103 == 1'h0;
  assign T_3156 = T_3145 & T_3155;
  assign T_3158 = T_3147 - 1'h1;
  assign T_3159 = T_3158[0:0];
  assign GEN_208 = T_3156 ? T_3159 : GEN_207;
  assign T_3161 = T_3147 > 1'h0;
  assign T_3162 = T_55 == 4'h6;
  assign T_3163 = T_175 >> T_186_up_idx;
  assign T_3164 = T_3163[0];
  assign T_3166 = T_3164 == 1'h0;
  assign T_3168 = T_59 | T_3166;
  assign T_3169 = T_3162 & T_3168;
  assign T_3172 = T_63 == 5'h1;
  assign T_3173 = T_63 == 5'h7;
  assign T_3174 = T_3172 | T_3173;
  assign T_3175 = T_63[3];
  assign T_3176 = T_63 == 5'h4;
  assign T_3177 = T_3175 | T_3176;
  assign T_3178 = T_3174 | T_3177;
  assign T_3179 = T_63 == 5'h3;
  assign T_3180 = T_3178 | T_3179;
  assign T_3181 = T_63 == 5'h6;
  assign T_3182 = T_3180 | T_3181;
  assign T_3185 = {T_63,1'h1};
  assign T_3216_addr_block = T_57;
  assign T_3216_client_xact_id = {{2'd0}, 1'h0};
  assign T_3216_addr_beat = {{2'd0}, 1'h0};
  assign T_3216_is_builtin_type = 1'h0;
  assign T_3216_a_type = {{2'd0}, T_3182};
  assign T_3216_union = {{6'd0}, T_3185};
  assign T_3216_data = {{63'd0}, 1'h0};
  assign GEN_11 = GEN_215;
  assign GEN_209 = GEN_444 == T_186_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_210 = GEN_465 == T_186_up_idx ? wmask_buffer_2 : GEN_209;
  assign GEN_211 = GEN_466 == T_186_up_idx ? wmask_buffer_3 : GEN_210;
  assign GEN_212 = 3'h4 == T_186_up_idx ? wmask_buffer_4 : GEN_211;
  assign GEN_213 = 3'h5 == T_186_up_idx ? wmask_buffer_5 : GEN_212;
  assign GEN_214 = 3'h6 == T_186_up_idx ? wmask_buffer_6 : GEN_213;
  assign GEN_215 = 3'h7 == T_186_up_idx ? wmask_buffer_7 : GEN_214;
  assign T_3281 = {T_63,1'h0};
  assign T_3282 = {T_65,T_67};
  assign T_3283 = {T_3282,T_3281};
  assign T_3285 = {T_67,T_63};
  assign T_3286 = {T_3285,1'h0};
  assign T_3288 = {GEN_11,1'h0};
  assign T_3300 = T_2111 ? 6'h2 : {{5'd0}, 1'h0};
  assign T_3302 = T_2113 ? 6'h0 : T_3300;
  assign T_3304 = T_2109 ? T_3283 : {{6'd0}, T_3302};
  assign T_3306 = T_2119 ? {{3'd0}, T_3288} : T_3304;
  assign T_3308 = T_2115 ? {{3'd0}, T_3288} : T_3306;
  assign T_3310 = T_2121 ? {{3'd0}, T_3286} : T_3308;
  assign T_3312 = T_2117 ? T_3283 : T_3310;
  assign T_3341_addr_block = T_57;
  assign T_3341_client_xact_id = {{2'd0}, 1'h0};
  assign T_3341_addr_beat = T_186_up_idx;
  assign T_3341_is_builtin_type = 1'h1;
  assign T_3341_a_type = T_99_a_type;
  assign T_3341_union = T_3312;
  assign T_3341_data = GEN_12;
  assign GEN_12 = GEN_222;
  assign GEN_216 = GEN_444 == T_186_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_217 = GEN_465 == T_186_up_idx ? data_buffer_2 : GEN_216;
  assign GEN_218 = GEN_466 == T_186_up_idx ? data_buffer_3 : GEN_217;
  assign GEN_219 = 3'h4 == T_186_up_idx ? data_buffer_4 : GEN_218;
  assign GEN_220 = 3'h5 == T_186_up_idx ? data_buffer_5 : GEN_219;
  assign GEN_221 = 3'h6 == T_186_up_idx ? data_buffer_6 : GEN_220;
  assign GEN_222 = 3'h7 == T_186_up_idx ? data_buffer_7 : GEN_221;
  assign T_3369_addr_block = T_3074 ? T_3216_addr_block : T_3341_addr_block;
  assign T_3369_client_xact_id = T_3074 ? T_3216_client_xact_id : T_3341_client_xact_id;
  assign T_3369_addr_beat = T_3074 ? T_3216_addr_beat : T_3341_addr_beat;
  assign T_3369_is_builtin_type = T_3074 ? T_3216_is_builtin_type : T_3341_is_builtin_type;
  assign T_3369_a_type = T_3074 ? T_3216_a_type : T_3341_a_type;
  assign T_3369_union = T_3074 ? T_3216_union : T_3341_union;
  assign T_3369_data = T_3074 ? T_3216_data : T_3341_data;
  assign T_3398 = T_3162 & T_186_up_done;
  assign GEN_223 = T_3398 ? 4'h7 : GEN_55;
  assign T_3408_0 = 3'h5;
  assign T_3408_1 = 3'h4;
  assign GEN_527 = {{1'd0}, T_3408_0};
  assign T_3410 = GEN_527 == io_outer_grant_bits_g_type;
  assign GEN_528 = {{1'd0}, T_3408_1};
  assign T_3411 = GEN_528 == io_outer_grant_bits_g_type;
  assign T_3414 = T_3410 | T_3411;
  assign T_3420_0 = 1'h0;
  assign GEN_529 = {{3'd0}, T_3420_0};
  assign T_3422 = GEN_529 == io_outer_grant_bits_g_type;
  assign T_3425 = io_outer_grant_bits_is_builtin_type ? T_3414 : T_3422;
  assign T_3426 = T_2405 & T_3425;
  assign GEN_13 = GEN_230;
  assign GEN_224 = GEN_444 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_225 = GEN_465 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_224;
  assign GEN_226 = GEN_466 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_225;
  assign GEN_227 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_226;
  assign GEN_228 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_227;
  assign GEN_229 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_228;
  assign GEN_230 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_229;
  assign T_3427 = GEN_13[0];
  assign GEN_14 = GEN_230;
  assign T_3428 = GEN_14[1];
  assign GEN_15 = GEN_230;
  assign T_3429 = GEN_15[2];
  assign GEN_16 = GEN_230;
  assign T_3430 = GEN_16[3];
  assign GEN_17 = GEN_230;
  assign T_3431 = GEN_17[4];
  assign GEN_18 = GEN_230;
  assign T_3432 = GEN_18[5];
  assign GEN_19 = GEN_230;
  assign T_3433 = GEN_19[6];
  assign GEN_20 = GEN_230;
  assign T_3434 = GEN_20[7];
  assign GEN_554 = {{7'd0}, T_3427};
  assign T_3436 = 8'h0 - GEN_554;
  assign T_3437 = T_3436[7:0];
  assign GEN_555 = {{7'd0}, T_3428};
  assign T_3439 = 8'h0 - GEN_555;
  assign T_3440 = T_3439[7:0];
  assign GEN_556 = {{7'd0}, T_3429};
  assign T_3442 = 8'h0 - GEN_556;
  assign T_3443 = T_3442[7:0];
  assign GEN_557 = {{7'd0}, T_3430};
  assign T_3445 = 8'h0 - GEN_557;
  assign T_3446 = T_3445[7:0];
  assign GEN_558 = {{7'd0}, T_3431};
  assign T_3448 = 8'h0 - GEN_558;
  assign T_3449 = T_3448[7:0];
  assign GEN_559 = {{7'd0}, T_3432};
  assign T_3451 = 8'h0 - GEN_559;
  assign T_3452 = T_3451[7:0];
  assign GEN_560 = {{7'd0}, T_3433};
  assign T_3454 = 8'h0 - GEN_560;
  assign T_3455 = T_3454[7:0];
  assign GEN_561 = {{7'd0}, T_3434};
  assign T_3457 = 8'h0 - GEN_561;
  assign T_3458 = T_3457[7:0];
  assign T_3464_0 = T_3437;
  assign T_3464_1 = T_3440;
  assign T_3464_2 = T_3443;
  assign T_3464_3 = T_3446;
  assign T_3464_4 = T_3449;
  assign T_3464_5 = T_3452;
  assign T_3464_6 = T_3455;
  assign T_3464_7 = T_3458;
  assign T_3466 = {T_3464_1,T_3464_0};
  assign T_3467 = {T_3464_3,T_3464_2};
  assign T_3468 = {T_3467,T_3466};
  assign T_3469 = {T_3464_5,T_3464_4};
  assign T_3470 = {T_3464_7,T_3464_6};
  assign T_3471 = {T_3470,T_3469};
  assign T_3472 = {T_3471,T_3468};
  assign T_3473 = ~ T_3472;
  assign T_3474 = T_3473 & io_outer_grant_bits_data;
  assign GEN_21 = GEN_286;
  assign GEN_280 = GEN_444 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_281 = GEN_465 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_280;
  assign GEN_282 = GEN_466 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_281;
  assign GEN_283 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_282;
  assign GEN_284 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_283;
  assign GEN_285 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_284;
  assign GEN_286 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_285;
  assign T_3475 = T_3472 & GEN_21;
  assign T_3476 = T_3474 | T_3475;
  assign GEN_22 = T_3476;
  assign GEN_287 = GEN_433 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_177;
  assign GEN_288 = GEN_444 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_178;
  assign GEN_289 = GEN_465 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_179;
  assign GEN_290 = GEN_466 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_180;
  assign GEN_291 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_181;
  assign GEN_292 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_182;
  assign GEN_293 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_183;
  assign GEN_294 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_22 : GEN_184;
  assign GEN_313 = T_3426 ? GEN_287 : GEN_177;
  assign GEN_314 = T_3426 ? GEN_288 : GEN_178;
  assign GEN_315 = T_3426 ? GEN_289 : GEN_179;
  assign GEN_316 = T_3426 ? GEN_290 : GEN_180;
  assign GEN_317 = T_3426 ? GEN_291 : GEN_181;
  assign GEN_318 = T_3426 ? GEN_292 : GEN_182;
  assign GEN_319 = T_3426 ? GEN_293 : GEN_183;
  assign GEN_320 = T_3426 ? GEN_294 : GEN_184;
  assign T_3477 = T_221 | T_186_pending;
  assign T_3478 = T_3477 | T_210_pending;
  assign T_3489 = T_2325 == 1'h0;
  assign T_3491 = T_2321 & T_3489;
  assign T_3499_0 = 3'h5;
  assign GEN_570 = {{1'd0}, T_3499_0};
  assign T_3501 = GEN_570 == io_inner_grant_bits_g_type;
  assign T_3509_0 = 2'h0;
  assign T_3509_1 = 2'h1;
  assign GEN_571 = {{2'd0}, T_3509_0};
  assign T_3511 = GEN_571 == io_inner_grant_bits_g_type;
  assign GEN_572 = {{2'd0}, T_3509_1};
  assign T_3512 = GEN_572 == io_inner_grant_bits_g_type;
  assign T_3515 = T_3511 | T_3512;
  assign T_3516 = io_inner_grant_bits_is_builtin_type ? T_3501 : T_3515;
  assign T_3518 = T_3491 & T_3516;
  assign T_3522 = T_3520 == 3'h7;
  assign T_3524 = T_3520 + GEN_444;
  assign T_3525 = T_3524[2:0];
  assign GEN_321 = T_3518 ? T_3525 : T_3520;
  assign T_3526 = T_3518 & T_3522;
  assign T_3527 = T_3516 ? T_3520 : {{2'd0}, 1'h0};
  assign T_3528 = T_3516 ? T_3526 : T_3491;
  assign T_3529 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3547 = T_3529 == 1'h0;
  assign T_3548 = T_3528 & T_3547;
  assign T_3550 = T_3545 + 1'h1;
  assign T_3551 = T_3550[0:0];
  assign GEN_323 = T_3548 ? T_3551 : T_3545;
  assign T_3553 = T_3528 == 1'h0;
  assign T_3554 = T_3529 & T_3553;
  assign T_3556 = T_3545 - 1'h1;
  assign T_3557 = T_3556[0:0];
  assign GEN_324 = T_3554 ? T_3557 : GEN_323;
  assign T_3559 = T_3545 > 1'h0;
  assign T_3564 = T_1885 == 1'h0;
  assign T_3573_0 = 3'h5;
  assign T_3573_1 = 3'h4;
  assign GEN_575 = {{1'd0}, T_3573_0};
  assign T_3575 = GEN_575 == io_inner_grant_bits_g_type;
  assign GEN_576 = {{1'd0}, T_3573_1};
  assign T_3576 = GEN_576 == io_inner_grant_bits_g_type;
  assign T_3579 = T_3575 | T_3576;
  assign T_3585_0 = 2'h0;
  assign T_3585_1 = 2'h1;
  assign GEN_577 = {{2'd0}, T_3585_0};
  assign T_3587 = GEN_577 == io_inner_grant_bits_g_type;
  assign GEN_578 = {{2'd0}, T_3585_1};
  assign T_3588 = GEN_578 == io_inner_grant_bits_g_type;
  assign T_3591 = T_3587 | T_3588;
  assign T_3592 = io_inner_grant_bits_is_builtin_type ? T_3579 : T_3591;
  assign T_3593 = T_2321 & T_3592;
  assign GEN_579 = {{7'd0}, T_3593};
  assign T_3595 = 8'h0 - GEN_579;
  assign T_3596 = T_3595[7:0];
  assign T_3597 = ~ T_3596;
  assign T_3599 = GEN_437 << io_inner_grant_bits_addr_beat;
  assign T_3600 = ~ T_3599;
  assign T_3601 = T_3597 | T_3600;
  assign T_3602 = T_177 & T_3601;
  assign T_3610_0 = 3'h0;
  assign T_3610_1 = 3'h1;
  assign T_3610_2 = 3'h2;
  assign T_3612 = T_3610_0 == io_inner_release_bits_r_type;
  assign T_3613 = T_3610_1 == io_inner_release_bits_r_type;
  assign T_3614 = T_3610_2 == io_inner_release_bits_r_type;
  assign T_3617 = T_3612 | T_3613;
  assign T_3618 = T_3617 | T_3614;
  assign T_3619 = T_2228 & T_3618;
  assign GEN_581 = {{7'd0}, T_3619};
  assign T_3622 = 8'h0 - GEN_581;
  assign T_3623 = T_3622[7:0];
  assign T_3626 = T_3623 & T_2476;
  assign T_3627 = T_3602 | T_3626;
  assign T_3637_0 = 3'h5;
  assign T_3637_1 = 3'h4;
  assign GEN_583 = {{1'd0}, T_3637_0};
  assign T_3639 = GEN_583 == io_outer_grant_bits_g_type;
  assign GEN_584 = {{1'd0}, T_3637_1};
  assign T_3640 = GEN_584 == io_outer_grant_bits_g_type;
  assign T_3643 = T_3639 | T_3640;
  assign T_3649_0 = 1'h0;
  assign GEN_585 = {{3'd0}, T_3649_0};
  assign T_3651 = GEN_585 == io_outer_grant_bits_g_type;
  assign T_3654 = io_outer_grant_bits_is_builtin_type ? T_3643 : T_3651;
  assign T_3655 = T_2405 & T_3654;
  assign GEN_586 = {{7'd0}, T_3655};
  assign T_3658 = 8'h0 - GEN_586;
  assign T_3659 = T_3658[7:0];
  assign T_3661 = GEN_437 << io_outer_grant_bits_addr_beat;
  assign T_3662 = T_3659 & T_3661;
  assign T_3663 = T_3627 | T_3662;
  assign T_3664 = T_3663 | GEN_432;
  assign GEN_335 = T_3564 ? T_3664 : GEN_43;
  assign T_3666 = T_55 == 4'h1;
  assign T_3667 = T_1733 | T_3666;
  assign T_3670 = T_3667 | T_2075;
  assign T_3672 = T_3670 == 1'h0;
  assign T_3689 = 3'h6 == Queue_14_1_io_deq_bits_a_type;
  assign T_3690 = T_3689 ? 3'h1 : 3'h3;
  assign T_3691 = 3'h5 == Queue_14_1_io_deq_bits_a_type;
  assign T_3692 = T_3691 ? 3'h1 : T_3690;
  assign T_3693 = 3'h4 == Queue_14_1_io_deq_bits_a_type;
  assign T_3694 = T_3693 ? 3'h4 : T_3692;
  assign T_3695 = 3'h3 == Queue_14_1_io_deq_bits_a_type;
  assign T_3696 = T_3695 ? 3'h3 : T_3694;
  assign T_3697 = 3'h2 == Queue_14_1_io_deq_bits_a_type;
  assign T_3698 = T_3697 ? 3'h3 : T_3696;
  assign T_3699 = 3'h1 == Queue_14_1_io_deq_bits_a_type;
  assign T_3700 = T_3699 ? 3'h5 : T_3698;
  assign T_3701 = 3'h0 == Queue_14_1_io_deq_bits_a_type;
  assign T_3702 = T_3701 ? 3'h4 : T_3700;
  assign T_3703 = Queue_14_1_io_deq_bits_a_type == GEN_433;
  assign T_3708 = T_3703 ? 2'h0 : 2'h1;
  assign T_3709 = Queue_14_1_io_deq_bits_is_builtin_type ? T_3702 : {{1'd0}, T_3708};
  assign T_3741_addr_beat = Queue_14_1_io_deq_bits_addr_beat;
  assign T_3741_client_xact_id = Queue_14_1_io_deq_bits_client_xact_id;
  assign T_3741_manager_xact_id = 3'h4;
  assign T_3741_is_builtin_type = Queue_14_1_io_deq_bits_is_builtin_type;
  assign T_3741_g_type = {{1'd0}, T_3709};
  assign T_3741_data = GEN_23;
  assign T_3741_client_id = Queue_14_1_io_deq_bits_client_id;
  assign GEN_23 = GEN_342;
  assign GEN_336 = GEN_444 == T_155 ? data_buffer_1 : data_buffer_0;
  assign GEN_337 = GEN_465 == T_155 ? data_buffer_2 : GEN_336;
  assign GEN_338 = GEN_466 == T_155 ? data_buffer_3 : GEN_337;
  assign GEN_339 = 3'h4 == T_155 ? data_buffer_4 : GEN_338;
  assign GEN_340 = 3'h5 == T_155 ? data_buffer_5 : GEN_339;
  assign GEN_341 = 3'h6 == T_155 ? data_buffer_6 : GEN_340;
  assign GEN_342 = 3'h7 == T_155 ? data_buffer_7 : GEN_341;
  assign T_3780_0 = 3'h5;
  assign GEN_594 = {{1'd0}, T_3780_0};
  assign T_3782 = GEN_594 == io_inner_grant_bits_g_type;
  assign T_3790_0 = 2'h0;
  assign T_3790_1 = 2'h1;
  assign GEN_595 = {{2'd0}, T_3790_0};
  assign T_3792 = GEN_595 == io_inner_grant_bits_g_type;
  assign GEN_596 = {{2'd0}, T_3790_1};
  assign T_3793 = GEN_596 == io_inner_grant_bits_g_type;
  assign T_3796 = T_3792 | T_3793;
  assign T_3797 = io_inner_grant_bits_is_builtin_type ? T_3782 : T_3796;
  assign T_3799 = T_2321 & T_3797;
  assign T_3803 = T_3801 == 3'h7;
  assign T_3805 = T_3801 + GEN_444;
  assign T_3806 = T_3805[2:0];
  assign GEN_343 = T_3799 ? T_3806 : T_3801;
  assign T_3807 = T_3799 & T_3803;
  assign T_3808 = T_3797 ? T_3801 : Queue_14_1_io_deq_bits_addr_beat;
  assign T_3809 = T_3797 ? T_3807 : T_2321;
  assign T_3814 = T_2977 & T_153;
  assign T_3816 = T_3478 == 1'h0;
  assign T_3824_0 = 3'h5;
  assign T_3824_1 = 3'h4;
  assign GEN_598 = {{1'd0}, T_3824_0};
  assign T_3826 = GEN_598 == io_inner_grant_bits_g_type;
  assign GEN_599 = {{1'd0}, T_3824_1};
  assign T_3827 = GEN_599 == io_inner_grant_bits_g_type;
  assign T_3830 = T_3826 | T_3827;
  assign T_3836_0 = 2'h0;
  assign T_3836_1 = 2'h1;
  assign GEN_600 = {{2'd0}, T_3836_0};
  assign T_3838 = GEN_600 == io_inner_grant_bits_g_type;
  assign GEN_601 = {{2'd0}, T_3836_1};
  assign T_3839 = GEN_601 == io_inner_grant_bits_g_type;
  assign T_3842 = T_3838 | T_3839;
  assign T_3843 = io_inner_grant_bits_is_builtin_type ? T_3830 : T_3842;
  assign T_3844 = T_177 >> T_155;
  assign T_3845 = T_3844[0];
  assign T_3846 = T_3843 ? T_3845 : T_3672;
  assign T_3847 = T_3816 & T_3846;
  assign GEN_348 = T_3814 ? T_3847 : T_2537;
  assign GEN_349 = T_2414 ? T_157 : 1'h0;
  assign GEN_350 = T_2414 ? T_155 : T_2639_addr_beat;
  assign GEN_351 = T_2414 ? T_3741_client_xact_id : T_2639_client_xact_id;
  assign GEN_352 = T_2414 ? T_3741_manager_xact_id : T_2639_manager_xact_id;
  assign GEN_353 = T_2414 ? T_3741_is_builtin_type : T_2639_is_builtin_type;
  assign GEN_354 = T_2414 ? T_3741_g_type : T_2639_g_type;
  assign GEN_355 = T_2414 ? T_3741_data : T_2639_data;
  assign GEN_356 = T_2414 ? T_3741_client_id : T_2639_client_id;
  assign GEN_361 = T_2414 ? GEN_348 : T_2537;
  assign T_3854 = ~ io_incoherent_0;
  assign GEN_362 = T_1885 ? {{1'd0}, T_3854} : T_2207;
  assign T_3869_0 = 3'h3;
  assign T_3871 = T_3869_0 == T_99_a_type;
  assign T_3874 = T_99_is_builtin_type & T_3871;
  assign T_3875 = T_1887 & T_3874;
  assign T_3876 = T_3875 & T_153;
  assign T_3879 = T_3876 & T_1905;
  assign T_3881 = T_3879 & io_inner_acquire_valid;
  assign T_3882 = T_1885 | T_3881;
  assign T_3892_0 = 3'h2;
  assign T_3892_1 = 3'h3;
  assign T_3892_2 = 3'h4;
  assign T_3894 = T_3892_0 == io_inner_acquire_bits_a_type;
  assign T_3895 = T_3892_1 == io_inner_acquire_bits_a_type;
  assign T_3896 = T_3892_2 == io_inner_acquire_bits_a_type;
  assign T_3899 = T_3894 | T_3895;
  assign T_3900 = T_3899 | T_3896;
  assign T_3901 = io_inner_acquire_bits_is_builtin_type & T_3900;
  assign T_3902 = T_1734 & T_3901;
  assign T_3903 = T_3902 & T_3882;
  assign T_3905 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3906 = io_inner_acquire_bits_is_builtin_type & T_3905;
  assign T_3910 = 8'h0 - GEN_437;
  assign T_3911 = T_3910[7:0];
  assign T_3917_0 = T_3911;
  assign T_3925 = T_2034 | T_2031;
  assign T_3926 = io_inner_acquire_bits_union[8:1];
  assign T_3928 = T_3925 ? T_3926 : {{7'd0}, 1'h0};
  assign T_3929 = T_3906 ? T_3917_0 : T_3928;
  assign T_3930 = T_3929[0];
  assign T_3931 = T_3929[1];
  assign T_3932 = T_3929[2];
  assign T_3933 = T_3929[3];
  assign T_3934 = T_3929[4];
  assign T_3935 = T_3929[5];
  assign T_3936 = T_3929[6];
  assign T_3937 = T_3929[7];
  assign GEN_603 = {{7'd0}, T_3930};
  assign T_3939 = 8'h0 - GEN_603;
  assign T_3940 = T_3939[7:0];
  assign GEN_604 = {{7'd0}, T_3931};
  assign T_3942 = 8'h0 - GEN_604;
  assign T_3943 = T_3942[7:0];
  assign GEN_605 = {{7'd0}, T_3932};
  assign T_3945 = 8'h0 - GEN_605;
  assign T_3946 = T_3945[7:0];
  assign GEN_606 = {{7'd0}, T_3933};
  assign T_3948 = 8'h0 - GEN_606;
  assign T_3949 = T_3948[7:0];
  assign GEN_607 = {{7'd0}, T_3934};
  assign T_3951 = 8'h0 - GEN_607;
  assign T_3952 = T_3951[7:0];
  assign GEN_608 = {{7'd0}, T_3935};
  assign T_3954 = 8'h0 - GEN_608;
  assign T_3955 = T_3954[7:0];
  assign GEN_609 = {{7'd0}, T_3936};
  assign T_3957 = 8'h0 - GEN_609;
  assign T_3958 = T_3957[7:0];
  assign GEN_610 = {{7'd0}, T_3937};
  assign T_3960 = 8'h0 - GEN_610;
  assign T_3961 = T_3960[7:0];
  assign T_3967_0 = T_3940;
  assign T_3967_1 = T_3943;
  assign T_3967_2 = T_3946;
  assign T_3967_3 = T_3949;
  assign T_3967_4 = T_3952;
  assign T_3967_5 = T_3955;
  assign T_3967_6 = T_3958;
  assign T_3967_7 = T_3961;
  assign T_3969 = {T_3967_1,T_3967_0};
  assign T_3970 = {T_3967_3,T_3967_2};
  assign T_3971 = {T_3970,T_3969};
  assign T_3972 = {T_3967_5,T_3967_4};
  assign T_3973 = {T_3967_7,T_3967_6};
  assign T_3974 = {T_3973,T_3972};
  assign T_3975 = {T_3974,T_3971};
  assign T_3976 = ~ T_3975;
  assign GEN_24 = GEN_369;
  assign GEN_363 = GEN_444 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_364 = GEN_465 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_363;
  assign GEN_365 = GEN_466 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_364;
  assign GEN_366 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_365;
  assign GEN_367 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_366;
  assign GEN_368 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_367;
  assign GEN_369 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_368;
  assign T_3977 = T_3976 & GEN_24;
  assign T_3978 = T_3975 & io_inner_acquire_bits_data;
  assign T_3979 = T_3977 | T_3978;
  assign GEN_25 = T_3979;
  assign GEN_370 = GEN_433 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_313;
  assign GEN_371 = GEN_444 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_314;
  assign GEN_372 = GEN_465 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_315;
  assign GEN_373 = GEN_466 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_316;
  assign GEN_374 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_317;
  assign GEN_375 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_318;
  assign GEN_376 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_319;
  assign GEN_377 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_25 : GEN_320;
  assign T_3993_0 = T_3911;
  assign T_4005 = T_3906 ? T_3993_0 : T_3928;
  assign GEN_26 = GEN_384;
  assign GEN_378 = GEN_444 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_379 = GEN_465 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_378;
  assign GEN_380 = GEN_466 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_379;
  assign GEN_381 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_380;
  assign GEN_382 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_381;
  assign GEN_383 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_382;
  assign GEN_384 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_383;
  assign T_4006 = T_4005 | GEN_26;
  assign GEN_27 = T_4006;
  assign GEN_385 = GEN_433 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_0;
  assign GEN_386 = GEN_444 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_1;
  assign GEN_387 = GEN_465 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_2;
  assign GEN_388 = GEN_466 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_3;
  assign GEN_389 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_4;
  assign GEN_390 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_5;
  assign GEN_391 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_6;
  assign GEN_392 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : wmask_buffer_7;
  assign GEN_404 = T_3903 ? GEN_370 : GEN_313;
  assign GEN_405 = T_3903 ? GEN_371 : GEN_314;
  assign GEN_406 = T_3903 ? GEN_372 : GEN_315;
  assign GEN_407 = T_3903 ? GEN_373 : GEN_316;
  assign GEN_408 = T_3903 ? GEN_374 : GEN_317;
  assign GEN_409 = T_3903 ? GEN_375 : GEN_318;
  assign GEN_410 = T_3903 ? GEN_376 : GEN_319;
  assign GEN_411 = T_3903 ? GEN_377 : GEN_320;
  assign GEN_415 = T_3903 ? GEN_385 : wmask_buffer_0;
  assign GEN_416 = T_3903 ? GEN_386 : wmask_buffer_1;
  assign GEN_417 = T_3903 ? GEN_387 : wmask_buffer_2;
  assign GEN_418 = T_3903 ? GEN_388 : wmask_buffer_3;
  assign GEN_419 = T_3903 ? GEN_389 : wmask_buffer_4;
  assign GEN_420 = T_3903 ? GEN_390 : wmask_buffer_5;
  assign GEN_421 = T_3903 ? GEN_391 : wmask_buffer_6;
  assign GEN_422 = T_3903 ? GEN_392 : wmask_buffer_7;
  assign T_4009 = T_2075 | T_2533;
  assign T_4010 = T_4009 | T_144_pending;
  assign T_4011 = T_4010 | T_221;
  assign T_4012 = T_4011 | T_210_pending;
  assign T_4013 = T_4012 | T_186_pending;
  assign T_4014 = T_4013 | T_153;
  assign T_4015 = T_4014 | T_166_pending;
  assign T_4017 = T_4015 == 1'h0;
  assign T_4019 = T_2977 & T_44;
  assign GEN_423 = T_4019 ? 4'h0 : GEN_223;
  assign GEN_424 = T_4019 ? {{7'd0}, 1'h0} : GEN_415;
  assign GEN_425 = T_4019 ? {{7'd0}, 1'h0} : GEN_416;
  assign GEN_426 = T_4019 ? {{7'd0}, 1'h0} : GEN_417;
  assign GEN_427 = T_4019 ? {{7'd0}, 1'h0} : GEN_418;
  assign GEN_428 = T_4019 ? {{7'd0}, 1'h0} : GEN_419;
  assign GEN_429 = T_4019 ? {{7'd0}, 1'h0} : GEN_420;
  assign GEN_430 = T_4019 ? {{7'd0}, 1'h0} : GEN_421;
  assign GEN_431 = T_4019 ? {{7'd0}, 1'h0} : GEN_422;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_30 = {1{$random}};
  T_55 = GEN_30[3:0];
  GEN_31 = {1{$random}};
  T_57 = GEN_31[25:0];
  GEN_39 = {1{$random}};
  T_59 = GEN_39[0:0];
  GEN_40 = {1{$random}};
  T_61 = GEN_40[4:0];
  GEN_41 = {1{$random}};
  T_63 = GEN_41[4:0];
  GEN_45 = {1{$random}};
  T_65 = GEN_45[2:0];
  GEN_59 = {1{$random}};
  T_67 = GEN_59[2:0];
  GEN_60 = {1{$random}};
  T_129 = GEN_60[2:0];
  GEN_61 = {1{$random}};
  T_131 = GEN_61[0:0];
  GEN_62 = {1{$random}};
  T_133 = GEN_62[1:0];
  GEN_63 = {1{$random}};
  T_135 = GEN_63[7:0];
  GEN_64 = {1{$random}};
  T_175 = GEN_64[7:0];
  GEN_66 = {1{$random}};
  T_177 = GEN_66[7:0];
  GEN_67 = {1{$random}};
  T_195 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  T_199 = GEN_68[0:0];
  GEN_70 = {1{$random}};
  T_201 = GEN_70[7:0];
  GEN_71 = {2{$random}};
  data_buffer_0 = GEN_71[63:0];
  GEN_72 = {2{$random}};
  data_buffer_1 = GEN_72[63:0];
  GEN_73 = {2{$random}};
  data_buffer_2 = GEN_73[63:0];
  GEN_74 = {2{$random}};
  data_buffer_3 = GEN_74[63:0];
  GEN_78 = {2{$random}};
  data_buffer_4 = GEN_78[63:0];
  GEN_79 = {2{$random}};
  data_buffer_5 = GEN_79[63:0];
  GEN_80 = {2{$random}};
  data_buffer_6 = GEN_80[63:0];
  GEN_81 = {2{$random}};
  data_buffer_7 = GEN_81[63:0];
  GEN_82 = {1{$random}};
  wmask_buffer_0 = GEN_82[7:0];
  GEN_83 = {1{$random}};
  wmask_buffer_1 = GEN_83[7:0];
  GEN_85 = {1{$random}};
  wmask_buffer_2 = GEN_85[7:0];
  GEN_86 = {1{$random}};
  wmask_buffer_3 = GEN_86[7:0];
  GEN_87 = {1{$random}};
  wmask_buffer_4 = GEN_87[7:0];
  GEN_95 = {1{$random}};
  wmask_buffer_5 = GEN_95[7:0];
  GEN_96 = {1{$random}};
  wmask_buffer_6 = GEN_96[7:0];
  GEN_97 = {1{$random}};
  wmask_buffer_7 = GEN_97[7:0];
  GEN_98 = {1{$random}};
  T_2219 = GEN_98[2:0];
  GEN_99 = {1{$random}};
  T_2252 = GEN_99[2:0];
  GEN_100 = {1{$random}};
  T_2262 = GEN_100[0:0];
  GEN_101 = {1{$random}};
  T_2312 = GEN_101[2:0];
  GEN_102 = {1{$random}};
  T_2356 = GEN_102[2:0];
  GEN_103 = {1{$random}};
  T_2366 = GEN_103[0:0];
  GEN_104 = {1{$random}};
  T_2912 = GEN_104[2:0];
  GEN_105 = {1{$random}};
  T_2952 = GEN_105[2:0];
  GEN_106 = {1{$random}};
  T_2962 = GEN_106[0:0];
  GEN_107 = {1{$random}};
  T_3095 = GEN_107[2:0];
  GEN_108 = {1{$random}};
  T_3137 = GEN_108[2:0];
  GEN_109 = {1{$random}};
  T_3147 = GEN_109[0:0];
  GEN_110 = {1{$random}};
  T_3520 = GEN_110[2:0];
  GEN_111 = {1{$random}};
  T_3535 = GEN_111[2:0];
  GEN_112 = {1{$random}};
  T_3545 = GEN_112[0:0];
  GEN_113 = {1{$random}};
  T_3801 = GEN_113[2:0];
  GEN_114 = {1{$random}};
  GEN_28 = GEN_114[0:0];
  GEN_115 = {1{$random}};
  GEN_29 = GEN_115[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_55 <= 4'h0;
    end else begin
      if(T_4019) begin
        T_55 <= 4'h0;
      end else begin
        if(T_3398) begin
          T_55 <= 4'h7;
        end else begin
          if(T_2383) begin
            T_55 <= 4'h7;
          end else begin
            if(T_2283) begin
              if(T_2183) begin
                T_55 <= 4'h6;
              end else begin
                T_55 <= 4'h7;
              end
            end else begin
              if(T_1885) begin
                T_55 <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_57 <= 26'h0;
    end else begin
      if(T_2383) begin
        T_57 <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1885) begin
          T_57 <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_59 <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_61 <= T_2028;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        if(T_2035) begin
          T_63 <= 5'h1;
        end else begin
          T_63 <= T_2036;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_65 <= T_2038;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1885) begin
        T_67 <= T_2039;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_129 <= io_inner_release_bits_r_type;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_131 <= io_inner_release_bits_client_id;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2228) begin
        if(T_2438) begin
          T_133 <= io_inner_release_bits_client_xact_id;
        end
      end
    end
    if(reset) begin
      T_135 <= 8'h0;
    end else begin
      if(T_2228) begin
        if(T_2489) begin
          T_135 <= T_2514;
        end else begin
          if(T_2438) begin
            if(T_2453) begin
              T_135 <= T_2478;
            end else begin
              T_135 <= {{7'd0}, 1'h0};
            end
          end
        end
      end
    end
    if(reset) begin
      T_175 <= 8'h0;
    end else begin
      if(T_1885) begin
        if(T_2034) begin
          T_175 <= T_2070;
        end else begin
          T_175 <= {{7'd0}, 1'h0};
        end
      end else begin
        if(T_1962) begin
          T_175 <= T_2020;
        end
      end
    end
    if(reset) begin
      T_177 <= 8'h0;
    end else begin
      if(T_3564) begin
        T_177 <= T_3664;
      end else begin
        if(T_1885) begin
          T_177 <= {{7'd0}, 1'h0};
        end
      end
    end
    if(1'h0) begin
    end else begin
      T_195 <= GEN_362[0];
    end
    if(reset) begin
      T_199 <= 1'h0;
    end else begin
      if(T_2833) begin
        T_199 <= 1'h0;
      end
    end
    if(reset) begin
      T_201 <= 8'h0;
    end else begin
      if(T_2832) begin
        T_201 <= T_2883;
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1817_0;
    end else begin
      if(T_3903) begin
        if(GEN_433 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_433 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_433 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_433 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_433 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_433 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_433 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1817_1;
    end else begin
      if(T_3903) begin
        if(GEN_444 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_444 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_444 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_444 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_444 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_444 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_444 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1817_2;
    end else begin
      if(T_3903) begin
        if(GEN_465 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_465 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_465 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_465 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_465 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_465 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_465 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1817_3;
    end else begin
      if(T_3903) begin
        if(GEN_466 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(GEN_466 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(GEN_466 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(GEN_466 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(GEN_466 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(GEN_466 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(GEN_466 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1817_4;
    end else begin
      if(T_3903) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1817_5;
    end else begin
      if(T_3903) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1817_6;
    end else begin
      if(T_3903) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1817_7;
    end else begin
      if(T_3903) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_25;
        end else begin
          if(T_3426) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_22;
            end else begin
              if(T_2725) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2725) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3426) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_22;
          end else begin
            if(T_2725) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2725) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1835_0;
    end else begin
      if(T_4019) begin
        wmask_buffer_0 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_433 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1835_1;
    end else begin
      if(T_4019) begin
        wmask_buffer_1 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_444 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1835_2;
    end else begin
      if(T_4019) begin
        wmask_buffer_2 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_465 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1835_3;
    end else begin
      if(T_4019) begin
        wmask_buffer_3 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(GEN_466 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1835_4;
    end else begin
      if(T_4019) begin
        wmask_buffer_4 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1835_5;
    end else begin
      if(T_4019) begin
        wmask_buffer_5 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1835_6;
    end else begin
      if(T_4019) begin
        wmask_buffer_6 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1835_7;
    end else begin
      if(T_4019) begin
        wmask_buffer_7 <= {{7'd0}, 1'h0};
      end else begin
        if(T_3903) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_27;
          end
        end
      end
    end
    if(reset) begin
      T_2219 <= 3'h0;
    end
    if(reset) begin
      T_2252 <= 3'h0;
    end else begin
      if(T_2250) begin
        T_2252 <= T_2257;
      end
    end
    if(reset) begin
      T_2262 <= 1'h0;
    end else begin
      if(T_2271) begin
        T_2262 <= T_2274;
      end else begin
        if(T_2265) begin
          T_2262 <= T_2268;
        end
      end
    end
    if(reset) begin
      T_2312 <= 3'h0;
    end else begin
      if(T_2310) begin
        T_2312 <= T_2317;
      end
    end
    if(reset) begin
      T_2356 <= 3'h0;
    end else begin
      if(T_2354) begin
        T_2356 <= T_2361;
      end
    end
    if(reset) begin
      T_2366 <= 1'h0;
    end else begin
      if(T_2375) begin
        T_2366 <= T_2378;
      end else begin
        if(T_2369) begin
          T_2366 <= T_2372;
        end
      end
    end
    if(reset) begin
      T_2912 <= 3'h0;
    end else begin
      if(T_2910) begin
        T_2912 <= T_2917;
      end
    end
    if(reset) begin
      T_2952 <= 3'h0;
    end else begin
      if(T_2950) begin
        T_2952 <= T_2957;
      end
    end
    if(reset) begin
      T_2962 <= 1'h0;
    end else begin
      if(T_2971) begin
        T_2962 <= T_2974;
      end else begin
        if(T_2965) begin
          T_2962 <= T_2968;
        end
      end
    end
    if(reset) begin
      T_3095 <= 3'h0;
    end else begin
      if(T_3093) begin
        T_3095 <= T_3100;
      end
    end
    if(reset) begin
      T_3137 <= 3'h0;
    end else begin
      if(T_3135) begin
        T_3137 <= T_3142;
      end
    end
    if(reset) begin
      T_3147 <= 1'h0;
    end else begin
      if(T_3156) begin
        T_3147 <= T_3159;
      end else begin
        if(T_3150) begin
          T_3147 <= T_3153;
        end
      end
    end
    if(reset) begin
      T_3520 <= 3'h0;
    end else begin
      if(T_3518) begin
        T_3520 <= T_3525;
      end
    end
    if(reset) begin
      T_3535 <= 3'h0;
    end
    if(reset) begin
      T_3545 <= 1'h0;
    end else begin
      if(T_3554) begin
        T_3545 <= T_3557;
      end else begin
        if(T_3548) begin
          T_3545 <= T_3551;
        end
      end
    end
    if(reset) begin
      T_3801 <= 3'h0;
    end else begin
      if(T_3799) begin
        T_3801 <= T_3806;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1778) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:95 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1778) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1778) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1792) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:99 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1792) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1792) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1803) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1803) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1803) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module LockingRRArbiter_5(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [2:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [11:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [2:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [11:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [2:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_addr_beat,
  input   io_in_2_bits_is_builtin_type,
  input  [2:0] io_in_2_bits_a_type,
  input  [11:0] io_in_2_bits_union,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [25:0] io_in_3_bits_addr_block,
  input  [2:0] io_in_3_bits_client_xact_id,
  input  [2:0] io_in_3_bits_addr_beat,
  input   io_in_3_bits_is_builtin_type,
  input  [2:0] io_in_3_bits_a_type,
  input  [11:0] io_in_3_bits_union,
  input  [63:0] io_in_3_bits_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [25:0] io_in_4_bits_addr_block,
  input  [2:0] io_in_4_bits_client_xact_id,
  input  [2:0] io_in_4_bits_addr_beat,
  input   io_in_4_bits_is_builtin_type,
  input  [2:0] io_in_4_bits_a_type,
  input  [11:0] io_in_4_bits_union,
  input  [63:0] io_in_4_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [2:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [11:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_52;
  wire  GEN_8;
  wire [2:0] GEN_53;
  wire  GEN_9;
  wire [2:0] GEN_54;
  wire  GEN_10;
  wire  GEN_11;
  wire [25:0] GEN_1;
  wire [25:0] GEN_12;
  wire [25:0] GEN_13;
  wire [25:0] GEN_14;
  wire [25:0] GEN_15;
  wire [2:0] GEN_2;
  wire [2:0] GEN_16;
  wire [2:0] GEN_17;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_3;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire  GEN_4;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire [2:0] GEN_5;
  wire [2:0] GEN_28;
  wire [2:0] GEN_29;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  wire [11:0] GEN_6;
  wire [11:0] GEN_32;
  wire [11:0] GEN_33;
  wire [11:0] GEN_34;
  wire [11:0] GEN_35;
  wire [63:0] GEN_7;
  wire [63:0] GEN_36;
  wire [63:0] GEN_37;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  reg [2:0] T_1114;
  reg [31:0] GEN_55;
  reg [2:0] T_1116;
  reg [31:0] GEN_56;
  wire [2:0] GEN_76;
  wire  T_1118;
  wire [2:0] T_1127_0;
  wire  T_1129;
  wire  T_1132;
  wire  T_1133;
  wire  T_1134;
  wire [3:0] T_1138;
  wire [2:0] T_1139;
  wire [2:0] GEN_40;
  wire [2:0] GEN_41;
  wire [2:0] GEN_42;
  reg [2:0] lastGrant;
  reg [31:0] GEN_57;
  wire [2:0] GEN_43;
  wire  T_1144;
  wire  T_1146;
  wire  T_1148;
  wire  T_1150;
  wire  T_1152;
  wire  T_1153;
  wire  T_1154;
  wire  T_1155;
  wire  T_1158;
  wire  T_1159;
  wire  T_1160;
  wire  T_1161;
  wire  T_1162;
  wire  T_1163;
  wire  T_1164;
  wire  T_1168;
  wire  T_1170;
  wire  T_1172;
  wire  T_1174;
  wire  T_1176;
  wire  T_1178;
  wire  T_1180;
  wire  T_1182;
  wire  T_1186;
  wire  T_1187;
  wire  T_1188;
  wire  T_1189;
  wire  T_1190;
  wire  T_1191;
  wire  T_1192;
  wire  T_1194;
  wire  T_1195;
  wire  T_1196;
  wire  T_1198;
  wire  T_1199;
  wire  T_1200;
  wire  T_1202;
  wire  T_1203;
  wire  T_1204;
  wire  T_1206;
  wire  T_1207;
  wire  T_1208;
  wire  T_1210;
  wire  T_1211;
  wire  T_1212;
  wire [2:0] GEN_44;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  wire [2:0] GEN_47;
  wire [2:0] GEN_48;
  wire [2:0] GEN_49;
  wire [2:0] GEN_50;
  wire [2:0] GEN_51;
  assign io_in_0_ready = T_1196;
  assign io_in_1_ready = T_1200;
  assign io_in_2_ready = T_1204;
  assign io_in_3_ready = T_1208;
  assign io_in_4_ready = T_1212;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_addr_beat = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_a_type = GEN_5;
  assign io_out_bits_union = GEN_6;
  assign io_out_bits_data = GEN_7;
  assign io_chosen = GEN_42;
  assign choice = GEN_51;
  assign GEN_0 = GEN_11;
  assign GEN_52 = {{2'd0}, 1'h1};
  assign GEN_8 = GEN_52 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_53 = {{1'd0}, 2'h2};
  assign GEN_9 = GEN_53 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_54 = {{1'd0}, 2'h3};
  assign GEN_10 = GEN_54 == io_chosen ? io_in_3_valid : GEN_9;
  assign GEN_11 = 3'h4 == io_chosen ? io_in_4_valid : GEN_10;
  assign GEN_1 = GEN_15;
  assign GEN_12 = GEN_52 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_13 = GEN_53 == io_chosen ? io_in_2_bits_addr_block : GEN_12;
  assign GEN_14 = GEN_54 == io_chosen ? io_in_3_bits_addr_block : GEN_13;
  assign GEN_15 = 3'h4 == io_chosen ? io_in_4_bits_addr_block : GEN_14;
  assign GEN_2 = GEN_19;
  assign GEN_16 = GEN_52 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_17 = GEN_53 == io_chosen ? io_in_2_bits_client_xact_id : GEN_16;
  assign GEN_18 = GEN_54 == io_chosen ? io_in_3_bits_client_xact_id : GEN_17;
  assign GEN_19 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_18;
  assign GEN_3 = GEN_23;
  assign GEN_20 = GEN_52 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_21 = GEN_53 == io_chosen ? io_in_2_bits_addr_beat : GEN_20;
  assign GEN_22 = GEN_54 == io_chosen ? io_in_3_bits_addr_beat : GEN_21;
  assign GEN_23 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_22;
  assign GEN_4 = GEN_27;
  assign GEN_24 = GEN_52 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_25 = GEN_53 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_24;
  assign GEN_26 = GEN_54 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_25;
  assign GEN_27 = 3'h4 == io_chosen ? io_in_4_bits_is_builtin_type : GEN_26;
  assign GEN_5 = GEN_31;
  assign GEN_28 = GEN_52 == io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_29 = GEN_53 == io_chosen ? io_in_2_bits_a_type : GEN_28;
  assign GEN_30 = GEN_54 == io_chosen ? io_in_3_bits_a_type : GEN_29;
  assign GEN_31 = 3'h4 == io_chosen ? io_in_4_bits_a_type : GEN_30;
  assign GEN_6 = GEN_35;
  assign GEN_32 = GEN_52 == io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_33 = GEN_53 == io_chosen ? io_in_2_bits_union : GEN_32;
  assign GEN_34 = GEN_54 == io_chosen ? io_in_3_bits_union : GEN_33;
  assign GEN_35 = 3'h4 == io_chosen ? io_in_4_bits_union : GEN_34;
  assign GEN_7 = GEN_39;
  assign GEN_36 = GEN_52 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_37 = GEN_53 == io_chosen ? io_in_2_bits_data : GEN_36;
  assign GEN_38 = GEN_54 == io_chosen ? io_in_3_bits_data : GEN_37;
  assign GEN_39 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_38;
  assign GEN_76 = {{2'd0}, 1'h0};
  assign T_1118 = T_1114 != GEN_76;
  assign T_1127_0 = 3'h3;
  assign T_1129 = T_1127_0 == io_out_bits_a_type;
  assign T_1132 = io_out_bits_is_builtin_type & T_1129;
  assign T_1133 = io_out_ready & io_out_valid;
  assign T_1134 = T_1133 & T_1132;
  assign T_1138 = T_1114 + GEN_52;
  assign T_1139 = T_1138[2:0];
  assign GEN_40 = T_1134 ? io_chosen : T_1116;
  assign GEN_41 = T_1134 ? T_1139 : T_1114;
  assign GEN_42 = T_1118 ? T_1116 : choice;
  assign GEN_43 = T_1133 ? io_chosen : lastGrant;
  assign T_1144 = GEN_52 > lastGrant;
  assign T_1146 = GEN_53 > lastGrant;
  assign T_1148 = GEN_54 > lastGrant;
  assign T_1150 = 3'h4 > lastGrant;
  assign T_1152 = io_in_1_valid & T_1144;
  assign T_1153 = io_in_2_valid & T_1146;
  assign T_1154 = io_in_3_valid & T_1148;
  assign T_1155 = io_in_4_valid & T_1150;
  assign T_1158 = T_1152 | T_1153;
  assign T_1159 = T_1158 | T_1154;
  assign T_1160 = T_1159 | T_1155;
  assign T_1161 = T_1160 | io_in_0_valid;
  assign T_1162 = T_1161 | io_in_1_valid;
  assign T_1163 = T_1162 | io_in_2_valid;
  assign T_1164 = T_1163 | io_in_3_valid;
  assign T_1168 = T_1152 == 1'h0;
  assign T_1170 = T_1158 == 1'h0;
  assign T_1172 = T_1159 == 1'h0;
  assign T_1174 = T_1160 == 1'h0;
  assign T_1176 = T_1161 == 1'h0;
  assign T_1178 = T_1162 == 1'h0;
  assign T_1180 = T_1163 == 1'h0;
  assign T_1182 = T_1164 == 1'h0;
  assign T_1186 = T_1144 | T_1176;
  assign T_1187 = T_1168 & T_1146;
  assign T_1188 = T_1187 | T_1178;
  assign T_1189 = T_1170 & T_1148;
  assign T_1190 = T_1189 | T_1180;
  assign T_1191 = T_1172 & T_1150;
  assign T_1192 = T_1191 | T_1182;
  assign T_1194 = T_1116 == GEN_76;
  assign T_1195 = T_1118 ? T_1194 : T_1174;
  assign T_1196 = T_1195 & io_out_ready;
  assign T_1198 = T_1116 == GEN_52;
  assign T_1199 = T_1118 ? T_1198 : T_1186;
  assign T_1200 = T_1199 & io_out_ready;
  assign T_1202 = T_1116 == GEN_53;
  assign T_1203 = T_1118 ? T_1202 : T_1188;
  assign T_1204 = T_1203 & io_out_ready;
  assign T_1206 = T_1116 == GEN_54;
  assign T_1207 = T_1118 ? T_1206 : T_1190;
  assign T_1208 = T_1207 & io_out_ready;
  assign T_1210 = T_1116 == 3'h4;
  assign T_1211 = T_1118 ? T_1210 : T_1192;
  assign T_1212 = T_1211 & io_out_ready;
  assign GEN_44 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_45 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_44;
  assign GEN_46 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_45;
  assign GEN_47 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_46;
  assign GEN_48 = T_1155 ? 3'h4 : GEN_47;
  assign GEN_49 = T_1154 ? {{1'd0}, 2'h3} : GEN_48;
  assign GEN_50 = T_1153 ? {{1'd0}, 2'h2} : GEN_49;
  assign GEN_51 = T_1152 ? {{2'd0}, 1'h1} : GEN_50;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_55 = {1{$random}};
  T_1114 = GEN_55[2:0];
  GEN_56 = {1{$random}};
  T_1116 = GEN_56[2:0];
  GEN_57 = {1{$random}};
  lastGrant = GEN_57[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1114 <= 3'h0;
    end else begin
      if(T_1134) begin
        T_1114 <= T_1139;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1134) begin
        T_1116 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1133) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module LockingRRArbiter_6(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [2:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [2:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [25:0] io_in_2_bits_addr_block,
  input  [2:0] io_in_2_bits_client_xact_id,
  input   io_in_2_bits_voluntary,
  input  [2:0] io_in_2_bits_r_type,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [25:0] io_in_3_bits_addr_block,
  input  [2:0] io_in_3_bits_client_xact_id,
  input   io_in_3_bits_voluntary,
  input  [2:0] io_in_3_bits_r_type,
  input  [63:0] io_in_3_bits_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_addr_beat,
  input  [25:0] io_in_4_bits_addr_block,
  input  [2:0] io_in_4_bits_client_xact_id,
  input   io_in_4_bits_voluntary,
  input  [2:0] io_in_4_bits_r_type,
  input  [63:0] io_in_4_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [2:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_47;
  wire  GEN_7;
  wire [2:0] GEN_48;
  wire  GEN_8;
  wire [2:0] GEN_49;
  wire  GEN_9;
  wire  GEN_10;
  wire [2:0] GEN_1;
  wire [2:0] GEN_11;
  wire [2:0] GEN_12;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [25:0] GEN_2;
  wire [25:0] GEN_15;
  wire [25:0] GEN_16;
  wire [25:0] GEN_17;
  wire [25:0] GEN_18;
  wire [2:0] GEN_3;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire  GEN_4;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire [2:0] GEN_5;
  wire [2:0] GEN_27;
  wire [2:0] GEN_28;
  wire [2:0] GEN_29;
  wire [2:0] GEN_30;
  wire [63:0] GEN_6;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  reg [2:0] T_1076;
  reg [31:0] GEN_50;
  reg [2:0] T_1078;
  reg [31:0] GEN_51;
  wire [2:0] GEN_68;
  wire  T_1080;
  wire [2:0] T_1087_0;
  wire [2:0] T_1087_1;
  wire [2:0] T_1087_2;
  wire  T_1089;
  wire  T_1090;
  wire  T_1091;
  wire  T_1094;
  wire  T_1095;
  wire  T_1097;
  wire  T_1098;
  wire [3:0] T_1102;
  wire [2:0] T_1103;
  wire [2:0] GEN_35;
  wire [2:0] GEN_36;
  wire [2:0] GEN_37;
  reg [2:0] lastGrant;
  reg [31:0] GEN_52;
  wire [2:0] GEN_38;
  wire  T_1108;
  wire  T_1110;
  wire  T_1112;
  wire  T_1114;
  wire  T_1116;
  wire  T_1117;
  wire  T_1118;
  wire  T_1119;
  wire  T_1122;
  wire  T_1123;
  wire  T_1124;
  wire  T_1125;
  wire  T_1126;
  wire  T_1127;
  wire  T_1128;
  wire  T_1132;
  wire  T_1134;
  wire  T_1136;
  wire  T_1138;
  wire  T_1140;
  wire  T_1142;
  wire  T_1144;
  wire  T_1146;
  wire  T_1150;
  wire  T_1151;
  wire  T_1152;
  wire  T_1153;
  wire  T_1154;
  wire  T_1155;
  wire  T_1156;
  wire  T_1158;
  wire  T_1159;
  wire  T_1160;
  wire  T_1162;
  wire  T_1163;
  wire  T_1164;
  wire  T_1166;
  wire  T_1167;
  wire  T_1168;
  wire  T_1170;
  wire  T_1171;
  wire  T_1172;
  wire  T_1174;
  wire  T_1175;
  wire  T_1176;
  wire [2:0] GEN_39;
  wire [2:0] GEN_40;
  wire [2:0] GEN_41;
  wire [2:0] GEN_42;
  wire [2:0] GEN_43;
  wire [2:0] GEN_44;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  assign io_in_0_ready = T_1160;
  assign io_in_1_ready = T_1164;
  assign io_in_2_ready = T_1168;
  assign io_in_3_ready = T_1172;
  assign io_in_4_ready = T_1176;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_addr_block = GEN_2;
  assign io_out_bits_client_xact_id = GEN_3;
  assign io_out_bits_voluntary = GEN_4;
  assign io_out_bits_r_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_37;
  assign choice = GEN_46;
  assign GEN_0 = GEN_10;
  assign GEN_47 = {{2'd0}, 1'h1};
  assign GEN_7 = GEN_47 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_48 = {{1'd0}, 2'h2};
  assign GEN_8 = GEN_48 == io_chosen ? io_in_2_valid : GEN_7;
  assign GEN_49 = {{1'd0}, 2'h3};
  assign GEN_9 = GEN_49 == io_chosen ? io_in_3_valid : GEN_8;
  assign GEN_10 = 3'h4 == io_chosen ? io_in_4_valid : GEN_9;
  assign GEN_1 = GEN_14;
  assign GEN_11 = GEN_47 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_12 = GEN_48 == io_chosen ? io_in_2_bits_addr_beat : GEN_11;
  assign GEN_13 = GEN_49 == io_chosen ? io_in_3_bits_addr_beat : GEN_12;
  assign GEN_14 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_13;
  assign GEN_2 = GEN_18;
  assign GEN_15 = GEN_47 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_16 = GEN_48 == io_chosen ? io_in_2_bits_addr_block : GEN_15;
  assign GEN_17 = GEN_49 == io_chosen ? io_in_3_bits_addr_block : GEN_16;
  assign GEN_18 = 3'h4 == io_chosen ? io_in_4_bits_addr_block : GEN_17;
  assign GEN_3 = GEN_22;
  assign GEN_19 = GEN_47 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_20 = GEN_48 == io_chosen ? io_in_2_bits_client_xact_id : GEN_19;
  assign GEN_21 = GEN_49 == io_chosen ? io_in_3_bits_client_xact_id : GEN_20;
  assign GEN_22 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_21;
  assign GEN_4 = GEN_26;
  assign GEN_23 = GEN_47 == io_chosen ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign GEN_24 = GEN_48 == io_chosen ? io_in_2_bits_voluntary : GEN_23;
  assign GEN_25 = GEN_49 == io_chosen ? io_in_3_bits_voluntary : GEN_24;
  assign GEN_26 = 3'h4 == io_chosen ? io_in_4_bits_voluntary : GEN_25;
  assign GEN_5 = GEN_30;
  assign GEN_27 = GEN_47 == io_chosen ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign GEN_28 = GEN_48 == io_chosen ? io_in_2_bits_r_type : GEN_27;
  assign GEN_29 = GEN_49 == io_chosen ? io_in_3_bits_r_type : GEN_28;
  assign GEN_30 = 3'h4 == io_chosen ? io_in_4_bits_r_type : GEN_29;
  assign GEN_6 = GEN_34;
  assign GEN_31 = GEN_47 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_32 = GEN_48 == io_chosen ? io_in_2_bits_data : GEN_31;
  assign GEN_33 = GEN_49 == io_chosen ? io_in_3_bits_data : GEN_32;
  assign GEN_34 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_33;
  assign GEN_68 = {{2'd0}, 1'h0};
  assign T_1080 = T_1076 != GEN_68;
  assign T_1087_0 = 3'h0;
  assign T_1087_1 = 3'h1;
  assign T_1087_2 = 3'h2;
  assign T_1089 = T_1087_0 == io_out_bits_r_type;
  assign T_1090 = T_1087_1 == io_out_bits_r_type;
  assign T_1091 = T_1087_2 == io_out_bits_r_type;
  assign T_1094 = T_1089 | T_1090;
  assign T_1095 = T_1094 | T_1091;
  assign T_1097 = io_out_ready & io_out_valid;
  assign T_1098 = T_1097 & T_1095;
  assign T_1102 = T_1076 + GEN_47;
  assign T_1103 = T_1102[2:0];
  assign GEN_35 = T_1098 ? io_chosen : T_1078;
  assign GEN_36 = T_1098 ? T_1103 : T_1076;
  assign GEN_37 = T_1080 ? T_1078 : choice;
  assign GEN_38 = T_1097 ? io_chosen : lastGrant;
  assign T_1108 = GEN_47 > lastGrant;
  assign T_1110 = GEN_48 > lastGrant;
  assign T_1112 = GEN_49 > lastGrant;
  assign T_1114 = 3'h4 > lastGrant;
  assign T_1116 = io_in_1_valid & T_1108;
  assign T_1117 = io_in_2_valid & T_1110;
  assign T_1118 = io_in_3_valid & T_1112;
  assign T_1119 = io_in_4_valid & T_1114;
  assign T_1122 = T_1116 | T_1117;
  assign T_1123 = T_1122 | T_1118;
  assign T_1124 = T_1123 | T_1119;
  assign T_1125 = T_1124 | io_in_0_valid;
  assign T_1126 = T_1125 | io_in_1_valid;
  assign T_1127 = T_1126 | io_in_2_valid;
  assign T_1128 = T_1127 | io_in_3_valid;
  assign T_1132 = T_1116 == 1'h0;
  assign T_1134 = T_1122 == 1'h0;
  assign T_1136 = T_1123 == 1'h0;
  assign T_1138 = T_1124 == 1'h0;
  assign T_1140 = T_1125 == 1'h0;
  assign T_1142 = T_1126 == 1'h0;
  assign T_1144 = T_1127 == 1'h0;
  assign T_1146 = T_1128 == 1'h0;
  assign T_1150 = T_1108 | T_1140;
  assign T_1151 = T_1132 & T_1110;
  assign T_1152 = T_1151 | T_1142;
  assign T_1153 = T_1134 & T_1112;
  assign T_1154 = T_1153 | T_1144;
  assign T_1155 = T_1136 & T_1114;
  assign T_1156 = T_1155 | T_1146;
  assign T_1158 = T_1078 == GEN_68;
  assign T_1159 = T_1080 ? T_1158 : T_1138;
  assign T_1160 = T_1159 & io_out_ready;
  assign T_1162 = T_1078 == GEN_47;
  assign T_1163 = T_1080 ? T_1162 : T_1150;
  assign T_1164 = T_1163 & io_out_ready;
  assign T_1166 = T_1078 == GEN_48;
  assign T_1167 = T_1080 ? T_1166 : T_1152;
  assign T_1168 = T_1167 & io_out_ready;
  assign T_1170 = T_1078 == GEN_49;
  assign T_1171 = T_1080 ? T_1170 : T_1154;
  assign T_1172 = T_1171 & io_out_ready;
  assign T_1174 = T_1078 == 3'h4;
  assign T_1175 = T_1080 ? T_1174 : T_1156;
  assign T_1176 = T_1175 & io_out_ready;
  assign GEN_39 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_40 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_39;
  assign GEN_41 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_40;
  assign GEN_42 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_41;
  assign GEN_43 = T_1119 ? 3'h4 : GEN_42;
  assign GEN_44 = T_1118 ? {{1'd0}, 2'h3} : GEN_43;
  assign GEN_45 = T_1117 ? {{1'd0}, 2'h2} : GEN_44;
  assign GEN_46 = T_1116 ? {{2'd0}, 1'h1} : GEN_45;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_50 = {1{$random}};
  T_1076 = GEN_50[2:0];
  GEN_51 = {1{$random}};
  T_1078 = GEN_51[2:0];
  GEN_52 = {1{$random}};
  lastGrant = GEN_52[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1076 <= 3'h0;
    end else begin
      if(T_1098) begin
        T_1076 <= T_1103;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1098) begin
        T_1078 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1097) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientTileLinkIOArbiter(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_probe_ready,
  output  io_in_0_probe_valid,
  output [25:0] io_in_0_probe_bits_addr_block,
  output [1:0] io_in_0_probe_bits_p_type,
  output  io_in_0_release_ready,
  input   io_in_0_release_valid,
  input  [2:0] io_in_0_release_bits_addr_beat,
  input  [25:0] io_in_0_release_bits_addr_block,
  input  [2:0] io_in_0_release_bits_client_xact_id,
  input   io_in_0_release_bits_voluntary,
  input  [2:0] io_in_0_release_bits_r_type,
  input  [63:0] io_in_0_release_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  output  io_in_0_grant_bits_manager_id,
  output  io_in_0_finish_ready,
  input   io_in_0_finish_valid,
  input   io_in_0_finish_bits_manager_xact_id,
  input   io_in_0_finish_bits_manager_id,
  output  io_in_1_acquire_ready,
  input   io_in_1_acquire_valid,
  input  [25:0] io_in_1_acquire_bits_addr_block,
  input  [2:0] io_in_1_acquire_bits_client_xact_id,
  input  [2:0] io_in_1_acquire_bits_addr_beat,
  input   io_in_1_acquire_bits_is_builtin_type,
  input  [2:0] io_in_1_acquire_bits_a_type,
  input  [11:0] io_in_1_acquire_bits_union,
  input  [63:0] io_in_1_acquire_bits_data,
  input   io_in_1_probe_ready,
  output  io_in_1_probe_valid,
  output [25:0] io_in_1_probe_bits_addr_block,
  output [1:0] io_in_1_probe_bits_p_type,
  output  io_in_1_release_ready,
  input   io_in_1_release_valid,
  input  [2:0] io_in_1_release_bits_addr_beat,
  input  [25:0] io_in_1_release_bits_addr_block,
  input  [2:0] io_in_1_release_bits_client_xact_id,
  input   io_in_1_release_bits_voluntary,
  input  [2:0] io_in_1_release_bits_r_type,
  input  [63:0] io_in_1_release_bits_data,
  input   io_in_1_grant_ready,
  output  io_in_1_grant_valid,
  output [2:0] io_in_1_grant_bits_addr_beat,
  output [2:0] io_in_1_grant_bits_client_xact_id,
  output  io_in_1_grant_bits_manager_xact_id,
  output  io_in_1_grant_bits_is_builtin_type,
  output [3:0] io_in_1_grant_bits_g_type,
  output [63:0] io_in_1_grant_bits_data,
  output  io_in_1_grant_bits_manager_id,
  output  io_in_1_finish_ready,
  input   io_in_1_finish_valid,
  input   io_in_1_finish_bits_manager_xact_id,
  input   io_in_1_finish_bits_manager_id,
  output  io_in_2_acquire_ready,
  input   io_in_2_acquire_valid,
  input  [25:0] io_in_2_acquire_bits_addr_block,
  input  [2:0] io_in_2_acquire_bits_client_xact_id,
  input  [2:0] io_in_2_acquire_bits_addr_beat,
  input   io_in_2_acquire_bits_is_builtin_type,
  input  [2:0] io_in_2_acquire_bits_a_type,
  input  [11:0] io_in_2_acquire_bits_union,
  input  [63:0] io_in_2_acquire_bits_data,
  input   io_in_2_probe_ready,
  output  io_in_2_probe_valid,
  output [25:0] io_in_2_probe_bits_addr_block,
  output [1:0] io_in_2_probe_bits_p_type,
  output  io_in_2_release_ready,
  input   io_in_2_release_valid,
  input  [2:0] io_in_2_release_bits_addr_beat,
  input  [25:0] io_in_2_release_bits_addr_block,
  input  [2:0] io_in_2_release_bits_client_xact_id,
  input   io_in_2_release_bits_voluntary,
  input  [2:0] io_in_2_release_bits_r_type,
  input  [63:0] io_in_2_release_bits_data,
  input   io_in_2_grant_ready,
  output  io_in_2_grant_valid,
  output [2:0] io_in_2_grant_bits_addr_beat,
  output [2:0] io_in_2_grant_bits_client_xact_id,
  output  io_in_2_grant_bits_manager_xact_id,
  output  io_in_2_grant_bits_is_builtin_type,
  output [3:0] io_in_2_grant_bits_g_type,
  output [63:0] io_in_2_grant_bits_data,
  output  io_in_2_grant_bits_manager_id,
  output  io_in_2_finish_ready,
  input   io_in_2_finish_valid,
  input   io_in_2_finish_bits_manager_xact_id,
  input   io_in_2_finish_bits_manager_id,
  output  io_in_3_acquire_ready,
  input   io_in_3_acquire_valid,
  input  [25:0] io_in_3_acquire_bits_addr_block,
  input  [2:0] io_in_3_acquire_bits_client_xact_id,
  input  [2:0] io_in_3_acquire_bits_addr_beat,
  input   io_in_3_acquire_bits_is_builtin_type,
  input  [2:0] io_in_3_acquire_bits_a_type,
  input  [11:0] io_in_3_acquire_bits_union,
  input  [63:0] io_in_3_acquire_bits_data,
  input   io_in_3_probe_ready,
  output  io_in_3_probe_valid,
  output [25:0] io_in_3_probe_bits_addr_block,
  output [1:0] io_in_3_probe_bits_p_type,
  output  io_in_3_release_ready,
  input   io_in_3_release_valid,
  input  [2:0] io_in_3_release_bits_addr_beat,
  input  [25:0] io_in_3_release_bits_addr_block,
  input  [2:0] io_in_3_release_bits_client_xact_id,
  input   io_in_3_release_bits_voluntary,
  input  [2:0] io_in_3_release_bits_r_type,
  input  [63:0] io_in_3_release_bits_data,
  input   io_in_3_grant_ready,
  output  io_in_3_grant_valid,
  output [2:0] io_in_3_grant_bits_addr_beat,
  output [2:0] io_in_3_grant_bits_client_xact_id,
  output  io_in_3_grant_bits_manager_xact_id,
  output  io_in_3_grant_bits_is_builtin_type,
  output [3:0] io_in_3_grant_bits_g_type,
  output [63:0] io_in_3_grant_bits_data,
  output  io_in_3_grant_bits_manager_id,
  output  io_in_3_finish_ready,
  input   io_in_3_finish_valid,
  input   io_in_3_finish_bits_manager_xact_id,
  input   io_in_3_finish_bits_manager_id,
  output  io_in_4_acquire_ready,
  input   io_in_4_acquire_valid,
  input  [25:0] io_in_4_acquire_bits_addr_block,
  input  [2:0] io_in_4_acquire_bits_client_xact_id,
  input  [2:0] io_in_4_acquire_bits_addr_beat,
  input   io_in_4_acquire_bits_is_builtin_type,
  input  [2:0] io_in_4_acquire_bits_a_type,
  input  [11:0] io_in_4_acquire_bits_union,
  input  [63:0] io_in_4_acquire_bits_data,
  input   io_in_4_probe_ready,
  output  io_in_4_probe_valid,
  output [25:0] io_in_4_probe_bits_addr_block,
  output [1:0] io_in_4_probe_bits_p_type,
  output  io_in_4_release_ready,
  input   io_in_4_release_valid,
  input  [2:0] io_in_4_release_bits_addr_beat,
  input  [25:0] io_in_4_release_bits_addr_block,
  input  [2:0] io_in_4_release_bits_client_xact_id,
  input   io_in_4_release_bits_voluntary,
  input  [2:0] io_in_4_release_bits_r_type,
  input  [63:0] io_in_4_release_bits_data,
  input   io_in_4_grant_ready,
  output  io_in_4_grant_valid,
  output [2:0] io_in_4_grant_bits_addr_beat,
  output [2:0] io_in_4_grant_bits_client_xact_id,
  output  io_in_4_grant_bits_manager_xact_id,
  output  io_in_4_grant_bits_is_builtin_type,
  output [3:0] io_in_4_grant_bits_g_type,
  output [63:0] io_in_4_grant_bits_data,
  output  io_in_4_grant_bits_manager_id,
  output  io_in_4_finish_ready,
  input   io_in_4_finish_valid,
  input   io_in_4_finish_bits_manager_xact_id,
  input   io_in_4_finish_bits_manager_id,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_probe_ready,
  input   io_out_probe_valid,
  input  [25:0] io_out_probe_bits_addr_block,
  input  [1:0] io_out_probe_bits_p_type,
  input   io_out_release_ready,
  output  io_out_release_valid,
  output [2:0] io_out_release_bits_addr_beat,
  output [25:0] io_out_release_bits_addr_block,
  output [2:0] io_out_release_bits_client_xact_id,
  output  io_out_release_bits_voluntary,
  output [2:0] io_out_release_bits_r_type,
  output [63:0] io_out_release_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data,
  input   io_out_grant_bits_manager_id,
  input   io_out_finish_ready,
  output  io_out_finish_valid,
  output  io_out_finish_bits_manager_xact_id,
  output  io_out_finish_bits_manager_id
);
  wire  LockingRRArbiter_5_1_clk;
  wire  LockingRRArbiter_5_1_reset;
  wire  LockingRRArbiter_5_1_io_in_0_ready;
  wire  LockingRRArbiter_5_1_io_in_0_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_0_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_0_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_0_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_0_bits_a_type;
  wire [11:0] LockingRRArbiter_5_1_io_in_0_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_0_bits_data;
  wire  LockingRRArbiter_5_1_io_in_1_ready;
  wire  LockingRRArbiter_5_1_io_in_1_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_1_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_1_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_1_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_1_bits_a_type;
  wire [11:0] LockingRRArbiter_5_1_io_in_1_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_1_bits_data;
  wire  LockingRRArbiter_5_1_io_in_2_ready;
  wire  LockingRRArbiter_5_1_io_in_2_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_2_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_2_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_2_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_2_bits_a_type;
  wire [11:0] LockingRRArbiter_5_1_io_in_2_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_2_bits_data;
  wire  LockingRRArbiter_5_1_io_in_3_ready;
  wire  LockingRRArbiter_5_1_io_in_3_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_3_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_3_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_3_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_3_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_3_bits_a_type;
  wire [11:0] LockingRRArbiter_5_1_io_in_3_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_3_bits_data;
  wire  LockingRRArbiter_5_1_io_in_4_ready;
  wire  LockingRRArbiter_5_1_io_in_4_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_4_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_4_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_4_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_4_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_4_bits_a_type;
  wire [11:0] LockingRRArbiter_5_1_io_in_4_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_4_bits_data;
  wire  LockingRRArbiter_5_1_io_out_ready;
  wire  LockingRRArbiter_5_1_io_out_valid;
  wire [25:0] LockingRRArbiter_5_1_io_out_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_out_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_out_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_out_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_out_bits_a_type;
  wire [11:0] LockingRRArbiter_5_1_io_out_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_out_bits_data;
  wire [2:0] LockingRRArbiter_5_1_io_chosen;
  wire [5:0] T_9040;
  wire [5:0] T_9042;
  wire [5:0] T_9044;
  wire [5:0] T_9046;
  wire [5:0] T_9048;
  wire  LockingRRArbiter_6_1_clk;
  wire  LockingRRArbiter_6_1_reset;
  wire  LockingRRArbiter_6_1_io_in_0_ready;
  wire  LockingRRArbiter_6_1_io_in_0_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_0_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_0_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_0_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_0_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_0_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_0_bits_data;
  wire  LockingRRArbiter_6_1_io_in_1_ready;
  wire  LockingRRArbiter_6_1_io_in_1_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_1_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_1_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_1_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_1_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_1_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_1_bits_data;
  wire  LockingRRArbiter_6_1_io_in_2_ready;
  wire  LockingRRArbiter_6_1_io_in_2_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_2_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_2_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_2_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_2_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_2_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_2_bits_data;
  wire  LockingRRArbiter_6_1_io_in_3_ready;
  wire  LockingRRArbiter_6_1_io_in_3_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_3_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_3_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_3_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_3_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_3_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_3_bits_data;
  wire  LockingRRArbiter_6_1_io_in_4_ready;
  wire  LockingRRArbiter_6_1_io_in_4_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_4_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_4_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_4_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_4_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_4_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_4_bits_data;
  wire  LockingRRArbiter_6_1_io_out_ready;
  wire  LockingRRArbiter_6_1_io_out_valid;
  wire [2:0] LockingRRArbiter_6_1_io_out_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_out_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_out_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_out_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_out_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_out_bits_data;
  wire [2:0] LockingRRArbiter_6_1_io_chosen;
  wire [5:0] T_9050;
  wire [5:0] T_9052;
  wire [5:0] T_9054;
  wire [5:0] T_9056;
  wire [5:0] T_9058;
  wire  T_9059;
  wire  T_9060;
  wire  T_9061;
  wire  T_9062;
  wire [2:0] GEN_10;
  wire  T_9067;
  wire  GEN_0;
  wire  GEN_1;
  wire [2:0] GEN_11;
  wire  T_9072;
  wire  GEN_2;
  wire  GEN_3;
  wire [2:0] GEN_12;
  wire  T_9077;
  wire  GEN_4;
  wire  GEN_5;
  wire [2:0] GEN_13;
  wire  T_9082;
  wire  GEN_6;
  wire  GEN_7;
  wire  T_9087;
  wire  GEN_8;
  wire  GEN_9;
  reg  GEN_14;
  reg [31:0] GEN_22;
  reg  GEN_15;
  reg [31:0] GEN_23;
  reg  GEN_16;
  reg [31:0] GEN_24;
  reg  GEN_17;
  reg [31:0] GEN_25;
  reg  GEN_18;
  reg [31:0] GEN_26;
  reg  GEN_19;
  reg [31:0] GEN_27;
  reg  GEN_20;
  reg [31:0] GEN_28;
  reg  GEN_21;
  reg [31:0] GEN_29;
  LockingRRArbiter_5 LockingRRArbiter_5_1 (
    .clk(LockingRRArbiter_5_1_clk),
    .reset(LockingRRArbiter_5_1_reset),
    .io_in_0_ready(LockingRRArbiter_5_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_5_1_io_in_0_valid),
    .io_in_0_bits_addr_block(LockingRRArbiter_5_1_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_5_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(LockingRRArbiter_5_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(LockingRRArbiter_5_1_io_in_0_bits_a_type),
    .io_in_0_bits_union(LockingRRArbiter_5_1_io_in_0_bits_union),
    .io_in_0_bits_data(LockingRRArbiter_5_1_io_in_0_bits_data),
    .io_in_1_ready(LockingRRArbiter_5_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_5_1_io_in_1_valid),
    .io_in_1_bits_addr_block(LockingRRArbiter_5_1_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_5_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(LockingRRArbiter_5_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(LockingRRArbiter_5_1_io_in_1_bits_a_type),
    .io_in_1_bits_union(LockingRRArbiter_5_1_io_in_1_bits_union),
    .io_in_1_bits_data(LockingRRArbiter_5_1_io_in_1_bits_data),
    .io_in_2_ready(LockingRRArbiter_5_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_5_1_io_in_2_valid),
    .io_in_2_bits_addr_block(LockingRRArbiter_5_1_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_5_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_addr_beat(LockingRRArbiter_5_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_a_type(LockingRRArbiter_5_1_io_in_2_bits_a_type),
    .io_in_2_bits_union(LockingRRArbiter_5_1_io_in_2_bits_union),
    .io_in_2_bits_data(LockingRRArbiter_5_1_io_in_2_bits_data),
    .io_in_3_ready(LockingRRArbiter_5_1_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_5_1_io_in_3_valid),
    .io_in_3_bits_addr_block(LockingRRArbiter_5_1_io_in_3_bits_addr_block),
    .io_in_3_bits_client_xact_id(LockingRRArbiter_5_1_io_in_3_bits_client_xact_id),
    .io_in_3_bits_addr_beat(LockingRRArbiter_5_1_io_in_3_bits_addr_beat),
    .io_in_3_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_a_type(LockingRRArbiter_5_1_io_in_3_bits_a_type),
    .io_in_3_bits_union(LockingRRArbiter_5_1_io_in_3_bits_union),
    .io_in_3_bits_data(LockingRRArbiter_5_1_io_in_3_bits_data),
    .io_in_4_ready(LockingRRArbiter_5_1_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_5_1_io_in_4_valid),
    .io_in_4_bits_addr_block(LockingRRArbiter_5_1_io_in_4_bits_addr_block),
    .io_in_4_bits_client_xact_id(LockingRRArbiter_5_1_io_in_4_bits_client_xact_id),
    .io_in_4_bits_addr_beat(LockingRRArbiter_5_1_io_in_4_bits_addr_beat),
    .io_in_4_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_4_bits_is_builtin_type),
    .io_in_4_bits_a_type(LockingRRArbiter_5_1_io_in_4_bits_a_type),
    .io_in_4_bits_union(LockingRRArbiter_5_1_io_in_4_bits_union),
    .io_in_4_bits_data(LockingRRArbiter_5_1_io_in_4_bits_data),
    .io_out_ready(LockingRRArbiter_5_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_5_1_io_out_valid),
    .io_out_bits_addr_block(LockingRRArbiter_5_1_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(LockingRRArbiter_5_1_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(LockingRRArbiter_5_1_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(LockingRRArbiter_5_1_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(LockingRRArbiter_5_1_io_out_bits_a_type),
    .io_out_bits_union(LockingRRArbiter_5_1_io_out_bits_union),
    .io_out_bits_data(LockingRRArbiter_5_1_io_out_bits_data),
    .io_chosen(LockingRRArbiter_5_1_io_chosen)
  );
  LockingRRArbiter_6 LockingRRArbiter_6_1 (
    .clk(LockingRRArbiter_6_1_clk),
    .reset(LockingRRArbiter_6_1_reset),
    .io_in_0_ready(LockingRRArbiter_6_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_6_1_io_in_0_valid),
    .io_in_0_bits_addr_beat(LockingRRArbiter_6_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(LockingRRArbiter_6_1_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_6_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(LockingRRArbiter_6_1_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(LockingRRArbiter_6_1_io_in_0_bits_r_type),
    .io_in_0_bits_data(LockingRRArbiter_6_1_io_in_0_bits_data),
    .io_in_1_ready(LockingRRArbiter_6_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_6_1_io_in_1_valid),
    .io_in_1_bits_addr_beat(LockingRRArbiter_6_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(LockingRRArbiter_6_1_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_6_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(LockingRRArbiter_6_1_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(LockingRRArbiter_6_1_io_in_1_bits_r_type),
    .io_in_1_bits_data(LockingRRArbiter_6_1_io_in_1_bits_data),
    .io_in_2_ready(LockingRRArbiter_6_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_6_1_io_in_2_valid),
    .io_in_2_bits_addr_beat(LockingRRArbiter_6_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_addr_block(LockingRRArbiter_6_1_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_6_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_voluntary(LockingRRArbiter_6_1_io_in_2_bits_voluntary),
    .io_in_2_bits_r_type(LockingRRArbiter_6_1_io_in_2_bits_r_type),
    .io_in_2_bits_data(LockingRRArbiter_6_1_io_in_2_bits_data),
    .io_in_3_ready(LockingRRArbiter_6_1_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_6_1_io_in_3_valid),
    .io_in_3_bits_addr_beat(LockingRRArbiter_6_1_io_in_3_bits_addr_beat),
    .io_in_3_bits_addr_block(LockingRRArbiter_6_1_io_in_3_bits_addr_block),
    .io_in_3_bits_client_xact_id(LockingRRArbiter_6_1_io_in_3_bits_client_xact_id),
    .io_in_3_bits_voluntary(LockingRRArbiter_6_1_io_in_3_bits_voluntary),
    .io_in_3_bits_r_type(LockingRRArbiter_6_1_io_in_3_bits_r_type),
    .io_in_3_bits_data(LockingRRArbiter_6_1_io_in_3_bits_data),
    .io_in_4_ready(LockingRRArbiter_6_1_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_6_1_io_in_4_valid),
    .io_in_4_bits_addr_beat(LockingRRArbiter_6_1_io_in_4_bits_addr_beat),
    .io_in_4_bits_addr_block(LockingRRArbiter_6_1_io_in_4_bits_addr_block),
    .io_in_4_bits_client_xact_id(LockingRRArbiter_6_1_io_in_4_bits_client_xact_id),
    .io_in_4_bits_voluntary(LockingRRArbiter_6_1_io_in_4_bits_voluntary),
    .io_in_4_bits_r_type(LockingRRArbiter_6_1_io_in_4_bits_r_type),
    .io_in_4_bits_data(LockingRRArbiter_6_1_io_in_4_bits_data),
    .io_out_ready(LockingRRArbiter_6_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_6_1_io_out_valid),
    .io_out_bits_addr_beat(LockingRRArbiter_6_1_io_out_bits_addr_beat),
    .io_out_bits_addr_block(LockingRRArbiter_6_1_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(LockingRRArbiter_6_1_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(LockingRRArbiter_6_1_io_out_bits_voluntary),
    .io_out_bits_r_type(LockingRRArbiter_6_1_io_out_bits_r_type),
    .io_out_bits_data(LockingRRArbiter_6_1_io_out_bits_data),
    .io_chosen(LockingRRArbiter_6_1_io_chosen)
  );
  assign io_in_0_acquire_ready = LockingRRArbiter_5_1_io_in_0_ready;
  assign io_in_0_probe_valid = io_out_probe_valid;
  assign io_in_0_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_0_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_0_release_ready = LockingRRArbiter_6_1_io_in_0_ready;
  assign io_in_0_grant_valid = GEN_0;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_0_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_0_finish_ready = GEN_14;
  assign io_in_1_acquire_ready = LockingRRArbiter_5_1_io_in_1_ready;
  assign io_in_1_probe_valid = io_out_probe_valid;
  assign io_in_1_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_1_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_1_release_ready = LockingRRArbiter_6_1_io_in_1_ready;
  assign io_in_1_grant_valid = GEN_2;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_1_finish_ready = GEN_15;
  assign io_in_2_acquire_ready = LockingRRArbiter_5_1_io_in_2_ready;
  assign io_in_2_probe_valid = io_out_probe_valid;
  assign io_in_2_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_2_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_2_release_ready = LockingRRArbiter_6_1_io_in_2_ready;
  assign io_in_2_grant_valid = GEN_4;
  assign io_in_2_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_2_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_2_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_2_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_2_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_2_grant_bits_data = io_out_grant_bits_data;
  assign io_in_2_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_2_finish_ready = GEN_16;
  assign io_in_3_acquire_ready = LockingRRArbiter_5_1_io_in_3_ready;
  assign io_in_3_probe_valid = io_out_probe_valid;
  assign io_in_3_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_3_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_3_release_ready = LockingRRArbiter_6_1_io_in_3_ready;
  assign io_in_3_grant_valid = GEN_6;
  assign io_in_3_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_3_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_3_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_3_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_3_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_3_grant_bits_data = io_out_grant_bits_data;
  assign io_in_3_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_3_finish_ready = GEN_17;
  assign io_in_4_acquire_ready = LockingRRArbiter_5_1_io_in_4_ready;
  assign io_in_4_probe_valid = io_out_probe_valid;
  assign io_in_4_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_4_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_4_release_ready = LockingRRArbiter_6_1_io_in_4_ready;
  assign io_in_4_grant_valid = GEN_8;
  assign io_in_4_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_4_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_4_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_4_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_4_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_4_grant_bits_data = io_out_grant_bits_data;
  assign io_in_4_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_4_finish_ready = GEN_18;
  assign io_out_acquire_valid = LockingRRArbiter_5_1_io_out_valid;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_5_1_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_5_1_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_5_1_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_5_1_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_5_1_io_out_bits_a_type;
  assign io_out_acquire_bits_union = LockingRRArbiter_5_1_io_out_bits_union;
  assign io_out_acquire_bits_data = LockingRRArbiter_5_1_io_out_bits_data;
  assign io_out_probe_ready = T_9062;
  assign io_out_release_valid = LockingRRArbiter_6_1_io_out_valid;
  assign io_out_release_bits_addr_beat = LockingRRArbiter_6_1_io_out_bits_addr_beat;
  assign io_out_release_bits_addr_block = LockingRRArbiter_6_1_io_out_bits_addr_block;
  assign io_out_release_bits_client_xact_id = LockingRRArbiter_6_1_io_out_bits_client_xact_id;
  assign io_out_release_bits_voluntary = LockingRRArbiter_6_1_io_out_bits_voluntary;
  assign io_out_release_bits_r_type = LockingRRArbiter_6_1_io_out_bits_r_type;
  assign io_out_release_bits_data = LockingRRArbiter_6_1_io_out_bits_data;
  assign io_out_grant_ready = GEN_9;
  assign io_out_finish_valid = GEN_19;
  assign io_out_finish_bits_manager_xact_id = GEN_20;
  assign io_out_finish_bits_manager_id = GEN_21;
  assign LockingRRArbiter_5_1_clk = clk;
  assign LockingRRArbiter_5_1_reset = reset;
  assign LockingRRArbiter_5_1_io_in_0_valid = io_in_0_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_0_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_0_bits_client_xact_id = T_9040[2:0];
  assign LockingRRArbiter_5_1_io_in_0_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_0_bits_a_type = io_in_0_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_0_bits_union = io_in_0_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_0_bits_data = io_in_0_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_1_valid = io_in_1_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_1_bits_addr_block = io_in_1_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_1_bits_client_xact_id = T_9042[2:0];
  assign LockingRRArbiter_5_1_io_in_1_bits_addr_beat = io_in_1_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type = io_in_1_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_1_bits_a_type = io_in_1_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_1_bits_union = io_in_1_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_1_bits_data = io_in_1_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_2_valid = io_in_2_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_2_bits_addr_block = io_in_2_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_2_bits_client_xact_id = T_9044[2:0];
  assign LockingRRArbiter_5_1_io_in_2_bits_addr_beat = io_in_2_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type = io_in_2_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_2_bits_a_type = io_in_2_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_2_bits_union = io_in_2_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_2_bits_data = io_in_2_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_3_valid = io_in_3_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_3_bits_addr_block = io_in_3_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_3_bits_client_xact_id = T_9046[2:0];
  assign LockingRRArbiter_5_1_io_in_3_bits_addr_beat = io_in_3_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_3_bits_is_builtin_type = io_in_3_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_3_bits_a_type = io_in_3_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_3_bits_union = io_in_3_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_3_bits_data = io_in_3_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_4_valid = io_in_4_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_4_bits_addr_block = io_in_4_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_4_bits_client_xact_id = T_9048[2:0];
  assign LockingRRArbiter_5_1_io_in_4_bits_addr_beat = io_in_4_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_4_bits_is_builtin_type = io_in_4_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_4_bits_a_type = io_in_4_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_4_bits_union = io_in_4_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_4_bits_data = io_in_4_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_out_ready = io_out_acquire_ready;
  assign T_9040 = {io_in_0_acquire_bits_client_xact_id,3'h0};
  assign T_9042 = {io_in_1_acquire_bits_client_xact_id,3'h1};
  assign T_9044 = {io_in_2_acquire_bits_client_xact_id,3'h2};
  assign T_9046 = {io_in_3_acquire_bits_client_xact_id,3'h3};
  assign T_9048 = {io_in_4_acquire_bits_client_xact_id,3'h4};
  assign LockingRRArbiter_6_1_clk = clk;
  assign LockingRRArbiter_6_1_reset = reset;
  assign LockingRRArbiter_6_1_io_in_0_valid = io_in_0_release_valid;
  assign LockingRRArbiter_6_1_io_in_0_bits_addr_beat = io_in_0_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_0_bits_addr_block = io_in_0_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_0_bits_client_xact_id = T_9050[2:0];
  assign LockingRRArbiter_6_1_io_in_0_bits_voluntary = io_in_0_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_0_bits_r_type = io_in_0_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_0_bits_data = io_in_0_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_1_valid = io_in_1_release_valid;
  assign LockingRRArbiter_6_1_io_in_1_bits_addr_beat = io_in_1_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_1_bits_addr_block = io_in_1_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_1_bits_client_xact_id = T_9052[2:0];
  assign LockingRRArbiter_6_1_io_in_1_bits_voluntary = io_in_1_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_1_bits_r_type = io_in_1_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_1_bits_data = io_in_1_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_2_valid = io_in_2_release_valid;
  assign LockingRRArbiter_6_1_io_in_2_bits_addr_beat = io_in_2_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_2_bits_addr_block = io_in_2_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_2_bits_client_xact_id = T_9054[2:0];
  assign LockingRRArbiter_6_1_io_in_2_bits_voluntary = io_in_2_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_2_bits_r_type = io_in_2_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_2_bits_data = io_in_2_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_3_valid = io_in_3_release_valid;
  assign LockingRRArbiter_6_1_io_in_3_bits_addr_beat = io_in_3_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_3_bits_addr_block = io_in_3_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_3_bits_client_xact_id = T_9056[2:0];
  assign LockingRRArbiter_6_1_io_in_3_bits_voluntary = io_in_3_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_3_bits_r_type = io_in_3_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_3_bits_data = io_in_3_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_4_valid = io_in_4_release_valid;
  assign LockingRRArbiter_6_1_io_in_4_bits_addr_beat = io_in_4_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_4_bits_addr_block = io_in_4_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_4_bits_client_xact_id = T_9058[2:0];
  assign LockingRRArbiter_6_1_io_in_4_bits_voluntary = io_in_4_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_4_bits_r_type = io_in_4_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_4_bits_data = io_in_4_release_bits_data;
  assign LockingRRArbiter_6_1_io_out_ready = io_out_release_ready;
  assign T_9050 = {io_in_0_release_bits_client_xact_id,3'h0};
  assign T_9052 = {io_in_1_release_bits_client_xact_id,3'h1};
  assign T_9054 = {io_in_2_release_bits_client_xact_id,3'h2};
  assign T_9056 = {io_in_3_release_bits_client_xact_id,3'h3};
  assign T_9058 = {io_in_4_release_bits_client_xact_id,3'h4};
  assign T_9059 = io_in_0_probe_ready & io_in_1_probe_ready;
  assign T_9060 = T_9059 & io_in_2_probe_ready;
  assign T_9061 = T_9060 & io_in_3_probe_ready;
  assign T_9062 = T_9061 & io_in_4_probe_ready;
  assign GEN_10 = {{2'd0}, 1'h0};
  assign T_9067 = io_out_grant_bits_client_xact_id == GEN_10;
  assign GEN_0 = T_9067 ? io_out_grant_valid : 1'h0;
  assign GEN_1 = T_9067 ? io_in_0_grant_ready : 1'h0;
  assign GEN_11 = {{2'd0}, 1'h1};
  assign T_9072 = io_out_grant_bits_client_xact_id == GEN_11;
  assign GEN_2 = T_9072 ? io_out_grant_valid : 1'h0;
  assign GEN_3 = T_9072 ? io_in_1_grant_ready : GEN_1;
  assign GEN_12 = {{1'd0}, 2'h2};
  assign T_9077 = io_out_grant_bits_client_xact_id == GEN_12;
  assign GEN_4 = T_9077 ? io_out_grant_valid : 1'h0;
  assign GEN_5 = T_9077 ? io_in_2_grant_ready : GEN_3;
  assign GEN_13 = {{1'd0}, 2'h3};
  assign T_9082 = io_out_grant_bits_client_xact_id == GEN_13;
  assign GEN_6 = T_9082 ? io_out_grant_valid : 1'h0;
  assign GEN_7 = T_9082 ? io_in_3_grant_ready : GEN_5;
  assign T_9087 = io_out_grant_bits_client_xact_id == 3'h4;
  assign GEN_8 = T_9087 ? io_out_grant_valid : 1'h0;
  assign GEN_9 = T_9087 ? io_in_4_grant_ready : GEN_7;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_22 = {1{$random}};
  GEN_14 = GEN_22[0:0];
  GEN_23 = {1{$random}};
  GEN_15 = GEN_23[0:0];
  GEN_24 = {1{$random}};
  GEN_16 = GEN_24[0:0];
  GEN_25 = {1{$random}};
  GEN_17 = GEN_25[0:0];
  GEN_26 = {1{$random}};
  GEN_18 = GEN_26[0:0];
  GEN_27 = {1{$random}};
  GEN_19 = GEN_27[0:0];
  GEN_28 = {1{$random}};
  GEN_20 = GEN_28[0:0];
  GEN_29 = {1{$random}};
  GEN_21 = GEN_29[0:0];
  end
`endif
endmodule
module LockingRRArbiter_7(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_p_type,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_p_type,
  input   io_in_1_bits_client_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_p_type,
  input   io_in_2_bits_client_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [25:0] io_in_3_bits_addr_block,
  input  [1:0] io_in_3_bits_p_type,
  input   io_in_3_bits_client_id,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [25:0] io_in_4_bits_addr_block,
  input  [1:0] io_in_4_bits_p_type,
  input   io_in_4_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_p_type,
  output  io_out_bits_client_id,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_32;
  wire  GEN_4;
  wire [2:0] GEN_33;
  wire  GEN_5;
  wire [2:0] GEN_34;
  wire  GEN_6;
  wire  GEN_7;
  wire [25:0] GEN_1;
  wire [25:0] GEN_8;
  wire [25:0] GEN_9;
  wire [25:0] GEN_10;
  wire [25:0] GEN_11;
  wire [1:0] GEN_2;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire  GEN_3;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  reg [2:0] T_1076;
  reg [31:0] GEN_20;
  reg [2:0] T_1078;
  reg [31:0] GEN_21;
  wire [2:0] GEN_44;
  wire  T_1080;
  wire  T_1082;
  wire [2:0] GEN_22;
  reg [2:0] lastGrant;
  reg [31:0] GEN_35;
  wire [2:0] GEN_23;
  wire  T_1093;
  wire  T_1095;
  wire  T_1097;
  wire  T_1099;
  wire  T_1101;
  wire  T_1102;
  wire  T_1103;
  wire  T_1104;
  wire  T_1107;
  wire  T_1108;
  wire  T_1109;
  wire  T_1110;
  wire  T_1111;
  wire  T_1112;
  wire  T_1113;
  wire  T_1117;
  wire  T_1119;
  wire  T_1121;
  wire  T_1123;
  wire  T_1125;
  wire  T_1127;
  wire  T_1129;
  wire  T_1131;
  wire  T_1135;
  wire  T_1136;
  wire  T_1137;
  wire  T_1138;
  wire  T_1139;
  wire  T_1140;
  wire  T_1141;
  wire  T_1143;
  wire  T_1144;
  wire  T_1145;
  wire  T_1147;
  wire  T_1148;
  wire  T_1149;
  wire  T_1151;
  wire  T_1152;
  wire  T_1153;
  wire  T_1155;
  wire  T_1156;
  wire  T_1157;
  wire  T_1159;
  wire  T_1160;
  wire  T_1161;
  wire [2:0] GEN_24;
  wire [2:0] GEN_25;
  wire [2:0] GEN_26;
  wire [2:0] GEN_27;
  wire [2:0] GEN_28;
  wire [2:0] GEN_29;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  assign io_in_0_ready = T_1145;
  assign io_in_1_ready = T_1149;
  assign io_in_2_ready = T_1153;
  assign io_in_3_ready = T_1157;
  assign io_in_4_ready = T_1161;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_p_type = GEN_2;
  assign io_out_bits_client_id = GEN_3;
  assign io_chosen = GEN_22;
  assign choice = GEN_31;
  assign GEN_0 = GEN_7;
  assign GEN_32 = {{2'd0}, 1'h1};
  assign GEN_4 = GEN_32 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_33 = {{1'd0}, 2'h2};
  assign GEN_5 = GEN_33 == io_chosen ? io_in_2_valid : GEN_4;
  assign GEN_34 = {{1'd0}, 2'h3};
  assign GEN_6 = GEN_34 == io_chosen ? io_in_3_valid : GEN_5;
  assign GEN_7 = 3'h4 == io_chosen ? io_in_4_valid : GEN_6;
  assign GEN_1 = GEN_11;
  assign GEN_8 = GEN_32 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_9 = GEN_33 == io_chosen ? io_in_2_bits_addr_block : GEN_8;
  assign GEN_10 = GEN_34 == io_chosen ? io_in_3_bits_addr_block : GEN_9;
  assign GEN_11 = 3'h4 == io_chosen ? io_in_4_bits_addr_block : GEN_10;
  assign GEN_2 = GEN_15;
  assign GEN_12 = GEN_32 == io_chosen ? io_in_1_bits_p_type : io_in_0_bits_p_type;
  assign GEN_13 = GEN_33 == io_chosen ? io_in_2_bits_p_type : GEN_12;
  assign GEN_14 = GEN_34 == io_chosen ? io_in_3_bits_p_type : GEN_13;
  assign GEN_15 = 3'h4 == io_chosen ? io_in_4_bits_p_type : GEN_14;
  assign GEN_3 = GEN_19;
  assign GEN_16 = GEN_32 == io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_17 = GEN_33 == io_chosen ? io_in_2_bits_client_id : GEN_16;
  assign GEN_18 = GEN_34 == io_chosen ? io_in_3_bits_client_id : GEN_17;
  assign GEN_19 = 3'h4 == io_chosen ? io_in_4_bits_client_id : GEN_18;
  assign GEN_44 = {{2'd0}, 1'h0};
  assign T_1080 = T_1076 != GEN_44;
  assign T_1082 = io_out_ready & io_out_valid;
  assign GEN_22 = T_1080 ? T_1078 : choice;
  assign GEN_23 = T_1082 ? io_chosen : lastGrant;
  assign T_1093 = GEN_32 > lastGrant;
  assign T_1095 = GEN_33 > lastGrant;
  assign T_1097 = GEN_34 > lastGrant;
  assign T_1099 = 3'h4 > lastGrant;
  assign T_1101 = io_in_1_valid & T_1093;
  assign T_1102 = io_in_2_valid & T_1095;
  assign T_1103 = io_in_3_valid & T_1097;
  assign T_1104 = io_in_4_valid & T_1099;
  assign T_1107 = T_1101 | T_1102;
  assign T_1108 = T_1107 | T_1103;
  assign T_1109 = T_1108 | T_1104;
  assign T_1110 = T_1109 | io_in_0_valid;
  assign T_1111 = T_1110 | io_in_1_valid;
  assign T_1112 = T_1111 | io_in_2_valid;
  assign T_1113 = T_1112 | io_in_3_valid;
  assign T_1117 = T_1101 == 1'h0;
  assign T_1119 = T_1107 == 1'h0;
  assign T_1121 = T_1108 == 1'h0;
  assign T_1123 = T_1109 == 1'h0;
  assign T_1125 = T_1110 == 1'h0;
  assign T_1127 = T_1111 == 1'h0;
  assign T_1129 = T_1112 == 1'h0;
  assign T_1131 = T_1113 == 1'h0;
  assign T_1135 = T_1093 | T_1125;
  assign T_1136 = T_1117 & T_1095;
  assign T_1137 = T_1136 | T_1127;
  assign T_1138 = T_1119 & T_1097;
  assign T_1139 = T_1138 | T_1129;
  assign T_1140 = T_1121 & T_1099;
  assign T_1141 = T_1140 | T_1131;
  assign T_1143 = T_1078 == GEN_44;
  assign T_1144 = T_1080 ? T_1143 : T_1123;
  assign T_1145 = T_1144 & io_out_ready;
  assign T_1147 = T_1078 == GEN_32;
  assign T_1148 = T_1080 ? T_1147 : T_1135;
  assign T_1149 = T_1148 & io_out_ready;
  assign T_1151 = T_1078 == GEN_33;
  assign T_1152 = T_1080 ? T_1151 : T_1137;
  assign T_1153 = T_1152 & io_out_ready;
  assign T_1155 = T_1078 == GEN_34;
  assign T_1156 = T_1080 ? T_1155 : T_1139;
  assign T_1157 = T_1156 & io_out_ready;
  assign T_1159 = T_1078 == 3'h4;
  assign T_1160 = T_1080 ? T_1159 : T_1141;
  assign T_1161 = T_1160 & io_out_ready;
  assign GEN_24 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_25 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_24;
  assign GEN_26 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_25;
  assign GEN_27 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_26;
  assign GEN_28 = T_1104 ? 3'h4 : GEN_27;
  assign GEN_29 = T_1103 ? {{1'd0}, 2'h3} : GEN_28;
  assign GEN_30 = T_1102 ? {{1'd0}, 2'h2} : GEN_29;
  assign GEN_31 = T_1101 ? {{2'd0}, 1'h1} : GEN_30;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_20 = {1{$random}};
  T_1076 = GEN_20[2:0];
  GEN_21 = {1{$random}};
  T_1078 = GEN_21[2:0];
  GEN_35 = {1{$random}};
  lastGrant = GEN_35[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1076 <= 3'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(T_1082) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module LockingRRArbiter_8(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [1:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  input   io_in_2_bits_client_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [1:0] io_in_3_bits_client_xact_id,
  input  [2:0] io_in_3_bits_manager_xact_id,
  input   io_in_3_bits_is_builtin_type,
  input  [3:0] io_in_3_bits_g_type,
  input  [63:0] io_in_3_bits_data,
  input   io_in_3_bits_client_id,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_addr_beat,
  input  [1:0] io_in_4_bits_client_xact_id,
  input  [2:0] io_in_4_bits_manager_xact_id,
  input   io_in_4_bits_is_builtin_type,
  input  [3:0] io_in_4_bits_g_type,
  input  [63:0] io_in_4_bits_data,
  input   io_in_4_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_52;
  wire  GEN_8;
  wire [2:0] GEN_53;
  wire  GEN_9;
  wire [2:0] GEN_54;
  wire  GEN_10;
  wire  GEN_11;
  wire [2:0] GEN_1;
  wire [2:0] GEN_12;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire [1:0] GEN_2;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [1:0] GEN_19;
  wire [2:0] GEN_3;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire  GEN_4;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire [3:0] GEN_5;
  wire [3:0] GEN_28;
  wire [3:0] GEN_29;
  wire [3:0] GEN_30;
  wire [3:0] GEN_31;
  wire [63:0] GEN_6;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire  GEN_7;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  reg [2:0] T_1228;
  reg [31:0] GEN_55;
  reg [2:0] T_1230;
  reg [31:0] GEN_56;
  wire [2:0] GEN_76;
  wire  T_1232;
  wire [2:0] T_1240_0;
  wire [3:0] GEN_77;
  wire  T_1242;
  wire [1:0] T_1250_0;
  wire [1:0] T_1250_1;
  wire [3:0] GEN_78;
  wire  T_1252;
  wire [3:0] GEN_79;
  wire  T_1253;
  wire  T_1256;
  wire  T_1257;
  wire  T_1259;
  wire  T_1260;
  wire [3:0] T_1264;
  wire [2:0] T_1265;
  wire [2:0] GEN_40;
  wire [2:0] GEN_41;
  wire [2:0] GEN_42;
  reg [2:0] lastGrant;
  reg [31:0] GEN_57;
  wire [2:0] GEN_43;
  wire  T_1270;
  wire  T_1272;
  wire  T_1274;
  wire  T_1276;
  wire  T_1278;
  wire  T_1279;
  wire  T_1280;
  wire  T_1281;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  wire  T_1287;
  wire  T_1288;
  wire  T_1289;
  wire  T_1290;
  wire  T_1294;
  wire  T_1296;
  wire  T_1298;
  wire  T_1300;
  wire  T_1302;
  wire  T_1304;
  wire  T_1306;
  wire  T_1308;
  wire  T_1312;
  wire  T_1313;
  wire  T_1314;
  wire  T_1315;
  wire  T_1316;
  wire  T_1317;
  wire  T_1318;
  wire  T_1320;
  wire  T_1321;
  wire  T_1322;
  wire  T_1324;
  wire  T_1325;
  wire  T_1326;
  wire  T_1328;
  wire  T_1329;
  wire  T_1330;
  wire  T_1332;
  wire  T_1333;
  wire  T_1334;
  wire  T_1336;
  wire  T_1337;
  wire  T_1338;
  wire [2:0] GEN_44;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  wire [2:0] GEN_47;
  wire [2:0] GEN_48;
  wire [2:0] GEN_49;
  wire [2:0] GEN_50;
  wire [2:0] GEN_51;
  assign io_in_0_ready = T_1322;
  assign io_in_1_ready = T_1326;
  assign io_in_2_ready = T_1330;
  assign io_in_3_ready = T_1334;
  assign io_in_4_ready = T_1338;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_client_id = GEN_7;
  assign io_chosen = GEN_42;
  assign choice = GEN_51;
  assign GEN_0 = GEN_11;
  assign GEN_52 = {{2'd0}, 1'h1};
  assign GEN_8 = GEN_52 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_53 = {{1'd0}, 2'h2};
  assign GEN_9 = GEN_53 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_54 = {{1'd0}, 2'h3};
  assign GEN_10 = GEN_54 == io_chosen ? io_in_3_valid : GEN_9;
  assign GEN_11 = 3'h4 == io_chosen ? io_in_4_valid : GEN_10;
  assign GEN_1 = GEN_15;
  assign GEN_12 = GEN_52 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_13 = GEN_53 == io_chosen ? io_in_2_bits_addr_beat : GEN_12;
  assign GEN_14 = GEN_54 == io_chosen ? io_in_3_bits_addr_beat : GEN_13;
  assign GEN_15 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_14;
  assign GEN_2 = GEN_19;
  assign GEN_16 = GEN_52 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_17 = GEN_53 == io_chosen ? io_in_2_bits_client_xact_id : GEN_16;
  assign GEN_18 = GEN_54 == io_chosen ? io_in_3_bits_client_xact_id : GEN_17;
  assign GEN_19 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_18;
  assign GEN_3 = GEN_23;
  assign GEN_20 = GEN_52 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_21 = GEN_53 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_20;
  assign GEN_22 = GEN_54 == io_chosen ? io_in_3_bits_manager_xact_id : GEN_21;
  assign GEN_23 = 3'h4 == io_chosen ? io_in_4_bits_manager_xact_id : GEN_22;
  assign GEN_4 = GEN_27;
  assign GEN_24 = GEN_52 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_25 = GEN_53 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_24;
  assign GEN_26 = GEN_54 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_25;
  assign GEN_27 = 3'h4 == io_chosen ? io_in_4_bits_is_builtin_type : GEN_26;
  assign GEN_5 = GEN_31;
  assign GEN_28 = GEN_52 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_29 = GEN_53 == io_chosen ? io_in_2_bits_g_type : GEN_28;
  assign GEN_30 = GEN_54 == io_chosen ? io_in_3_bits_g_type : GEN_29;
  assign GEN_31 = 3'h4 == io_chosen ? io_in_4_bits_g_type : GEN_30;
  assign GEN_6 = GEN_35;
  assign GEN_32 = GEN_52 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_33 = GEN_53 == io_chosen ? io_in_2_bits_data : GEN_32;
  assign GEN_34 = GEN_54 == io_chosen ? io_in_3_bits_data : GEN_33;
  assign GEN_35 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_34;
  assign GEN_7 = GEN_39;
  assign GEN_36 = GEN_52 == io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_37 = GEN_53 == io_chosen ? io_in_2_bits_client_id : GEN_36;
  assign GEN_38 = GEN_54 == io_chosen ? io_in_3_bits_client_id : GEN_37;
  assign GEN_39 = 3'h4 == io_chosen ? io_in_4_bits_client_id : GEN_38;
  assign GEN_76 = {{2'd0}, 1'h0};
  assign T_1232 = T_1228 != GEN_76;
  assign T_1240_0 = 3'h5;
  assign GEN_77 = {{1'd0}, T_1240_0};
  assign T_1242 = GEN_77 == io_out_bits_g_type;
  assign T_1250_0 = 2'h0;
  assign T_1250_1 = 2'h1;
  assign GEN_78 = {{2'd0}, T_1250_0};
  assign T_1252 = GEN_78 == io_out_bits_g_type;
  assign GEN_79 = {{2'd0}, T_1250_1};
  assign T_1253 = GEN_79 == io_out_bits_g_type;
  assign T_1256 = T_1252 | T_1253;
  assign T_1257 = io_out_bits_is_builtin_type ? T_1242 : T_1256;
  assign T_1259 = io_out_ready & io_out_valid;
  assign T_1260 = T_1259 & T_1257;
  assign T_1264 = T_1228 + GEN_52;
  assign T_1265 = T_1264[2:0];
  assign GEN_40 = T_1260 ? io_chosen : T_1230;
  assign GEN_41 = T_1260 ? T_1265 : T_1228;
  assign GEN_42 = T_1232 ? T_1230 : choice;
  assign GEN_43 = T_1259 ? io_chosen : lastGrant;
  assign T_1270 = GEN_52 > lastGrant;
  assign T_1272 = GEN_53 > lastGrant;
  assign T_1274 = GEN_54 > lastGrant;
  assign T_1276 = 3'h4 > lastGrant;
  assign T_1278 = io_in_1_valid & T_1270;
  assign T_1279 = io_in_2_valid & T_1272;
  assign T_1280 = io_in_3_valid & T_1274;
  assign T_1281 = io_in_4_valid & T_1276;
  assign T_1284 = T_1278 | T_1279;
  assign T_1285 = T_1284 | T_1280;
  assign T_1286 = T_1285 | T_1281;
  assign T_1287 = T_1286 | io_in_0_valid;
  assign T_1288 = T_1287 | io_in_1_valid;
  assign T_1289 = T_1288 | io_in_2_valid;
  assign T_1290 = T_1289 | io_in_3_valid;
  assign T_1294 = T_1278 == 1'h0;
  assign T_1296 = T_1284 == 1'h0;
  assign T_1298 = T_1285 == 1'h0;
  assign T_1300 = T_1286 == 1'h0;
  assign T_1302 = T_1287 == 1'h0;
  assign T_1304 = T_1288 == 1'h0;
  assign T_1306 = T_1289 == 1'h0;
  assign T_1308 = T_1290 == 1'h0;
  assign T_1312 = T_1270 | T_1302;
  assign T_1313 = T_1294 & T_1272;
  assign T_1314 = T_1313 | T_1304;
  assign T_1315 = T_1296 & T_1274;
  assign T_1316 = T_1315 | T_1306;
  assign T_1317 = T_1298 & T_1276;
  assign T_1318 = T_1317 | T_1308;
  assign T_1320 = T_1230 == GEN_76;
  assign T_1321 = T_1232 ? T_1320 : T_1300;
  assign T_1322 = T_1321 & io_out_ready;
  assign T_1324 = T_1230 == GEN_52;
  assign T_1325 = T_1232 ? T_1324 : T_1312;
  assign T_1326 = T_1325 & io_out_ready;
  assign T_1328 = T_1230 == GEN_53;
  assign T_1329 = T_1232 ? T_1328 : T_1314;
  assign T_1330 = T_1329 & io_out_ready;
  assign T_1332 = T_1230 == GEN_54;
  assign T_1333 = T_1232 ? T_1332 : T_1316;
  assign T_1334 = T_1333 & io_out_ready;
  assign T_1336 = T_1230 == 3'h4;
  assign T_1337 = T_1232 ? T_1336 : T_1318;
  assign T_1338 = T_1337 & io_out_ready;
  assign GEN_44 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_45 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_44;
  assign GEN_46 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_45;
  assign GEN_47 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_46;
  assign GEN_48 = T_1281 ? 3'h4 : GEN_47;
  assign GEN_49 = T_1280 ? {{1'd0}, 2'h3} : GEN_48;
  assign GEN_50 = T_1279 ? {{1'd0}, 2'h2} : GEN_49;
  assign GEN_51 = T_1278 ? {{2'd0}, 1'h1} : GEN_50;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_55 = {1{$random}};
  T_1228 = GEN_55[2:0];
  GEN_56 = {1{$random}};
  T_1230 = GEN_56[2:0];
  GEN_57 = {1{$random}};
  lastGrant = GEN_57[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1228 <= 3'h0;
    end else begin
      if(T_1260) begin
        T_1228 <= T_1265;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1260) begin
        T_1230 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1259) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module L2BroadcastHub(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_clk;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_reset;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_valid;
  wire [25:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_addr_block;
  wire [1:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_addr_beat;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_union;
  wire [63:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_data;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_client_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_valid;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_addr_beat;
  wire [1:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_manager_xact_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_g_type;
  wire [63:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_data;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_client_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_valid;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_bits_manager_xact_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_valid;
  wire [25:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_p_type;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_client_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_valid;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_addr_block;
  wire [1:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_client_xact_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_voluntary;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_r_type;
  wire [63:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_data;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_client_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_incoherent_0;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_valid;
  wire [25:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_addr_block;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_addr_beat;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_union;
  wire [63:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_data;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_valid;
  wire [25:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_bits_p_type;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_valid;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_addr_block;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_client_xact_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_voluntary;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_r_type;
  wire [63:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_data;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_valid;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_addr_beat;
  wire [2:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_client_xact_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_manager_xact_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_g_type;
  wire [63:0] BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_data;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_manager_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_ready;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_valid;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_bits_manager_xact_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_bits_manager_id;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_matches;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_can;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_should;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_matches;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_can;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_should;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_oprb_matches;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_oprb_can;
  wire  BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_oprb_should;
  wire  BufferedBroadcastAcquireTracker_4_clk;
  wire  BufferedBroadcastAcquireTracker_4_reset;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_acquire_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_acquire_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_addr_beat;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_union;
  wire [63:0] BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_data;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_grant_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_grant_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat;
  wire [1:0] BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_g_type;
  wire [63:0] BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_data;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_finish_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_finish_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_inner_finish_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_probe_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_probe_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_p_type;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_release_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_release_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_inner_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastAcquireTracker_4_io_inner_release_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_4_io_inner_release_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_release_bits_voluntary;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_inner_release_bits_r_type;
  wire [63:0] BufferedBroadcastAcquireTracker_4_io_inner_release_bits_data;
  wire  BufferedBroadcastAcquireTracker_4_io_inner_release_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_4_io_incoherent_0;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_acquire_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_acquire_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_union;
  wire [63:0] BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_data;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_probe_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_probe_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_4_io_outer_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_4_io_outer_probe_bits_p_type;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_release_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_release_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_outer_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastAcquireTracker_4_io_outer_release_bits_addr_block;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_outer_release_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_release_bits_voluntary;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_outer_release_bits_r_type;
  wire [63:0] BufferedBroadcastAcquireTracker_4_io_outer_release_bits_data;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_grant_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_grant_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_addr_beat;
  wire [2:0] BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_g_type;
  wire [63:0] BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_data;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_manager_id;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_finish_ready;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_finish_valid;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_finish_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_4_io_outer_finish_bits_manager_id;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_iacq_matches;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_iacq_can;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_iacq_should;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_irel_matches;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_irel_can;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_irel_should;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_oprb_matches;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_oprb_can;
  wire  BufferedBroadcastAcquireTracker_4_io_alloc_oprb_should;
  wire  BufferedBroadcastAcquireTracker_1_1_clk;
  wire  BufferedBroadcastAcquireTracker_1_1_reset;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_addr_beat;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_union;
  wire [63:0] BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_data;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_grant_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_grant_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_addr_beat;
  wire [1:0] BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_g_type;
  wire [63:0] BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_data;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_finish_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_finish_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_inner_finish_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_probe_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_probe_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_p_type;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_release_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_release_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_voluntary;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_r_type;
  wire [63:0] BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_data;
  wire  BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_incoherent_0;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_addr_block;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_addr_beat;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_union;
  wire [63:0] BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_data;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_probe_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_probe_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_1_1_io_outer_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_1_1_io_outer_probe_bits_p_type;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_release_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_release_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_addr_block;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_voluntary;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_r_type;
  wire [63:0] BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_data;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_grant_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_grant_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_addr_beat;
  wire [2:0] BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_g_type;
  wire [63:0] BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_data;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_manager_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_finish_ready;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_finish_valid;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_finish_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_outer_finish_bits_manager_id;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_matches;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_can;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_should;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_matches;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_can;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_should;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_oprb_matches;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_oprb_can;
  wire  BufferedBroadcastAcquireTracker_1_1_io_alloc_oprb_should;
  wire  BufferedBroadcastAcquireTracker_2_1_clk;
  wire  BufferedBroadcastAcquireTracker_2_1_reset;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_addr_beat;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_union;
  wire [63:0] BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_data;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_grant_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_grant_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_addr_beat;
  wire [1:0] BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_g_type;
  wire [63:0] BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_data;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_finish_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_finish_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_inner_finish_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_probe_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_probe_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_p_type;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_release_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_release_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_voluntary;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_r_type;
  wire [63:0] BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_data;
  wire  BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_incoherent_0;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_addr_block;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_addr_beat;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_union;
  wire [63:0] BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_data;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_probe_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_probe_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_2_1_io_outer_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_2_1_io_outer_probe_bits_p_type;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_release_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_release_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_addr_block;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_voluntary;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_r_type;
  wire [63:0] BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_data;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_grant_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_grant_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_addr_beat;
  wire [2:0] BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_g_type;
  wire [63:0] BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_data;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_manager_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_finish_ready;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_finish_valid;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_finish_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_outer_finish_bits_manager_id;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_matches;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_can;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_should;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_matches;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_can;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_should;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_oprb_matches;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_oprb_can;
  wire  BufferedBroadcastAcquireTracker_2_1_io_alloc_oprb_should;
  wire  BufferedBroadcastAcquireTracker_3_1_clk;
  wire  BufferedBroadcastAcquireTracker_3_1_reset;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_addr_beat;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_union;
  wire [63:0] BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_data;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_grant_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_grant_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_addr_beat;
  wire [1:0] BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_g_type;
  wire [63:0] BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_data;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_finish_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_finish_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_inner_finish_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_probe_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_probe_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_p_type;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_release_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_release_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_voluntary;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_r_type;
  wire [63:0] BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_data;
  wire  BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_client_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_incoherent_0;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_addr_block;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_addr_beat;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_a_type;
  wire [11:0] BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_union;
  wire [63:0] BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_data;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_probe_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_probe_valid;
  wire [25:0] BufferedBroadcastAcquireTracker_3_1_io_outer_probe_bits_addr_block;
  wire [1:0] BufferedBroadcastAcquireTracker_3_1_io_outer_probe_bits_p_type;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_release_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_release_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_addr_beat;
  wire [25:0] BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_addr_block;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_voluntary;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_r_type;
  wire [63:0] BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_data;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_grant_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_grant_valid;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_addr_beat;
  wire [2:0] BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_client_xact_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_g_type;
  wire [63:0] BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_data;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_manager_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_finish_ready;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_finish_valid;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_finish_bits_manager_xact_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_outer_finish_bits_manager_id;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_matches;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_can;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_should;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_matches;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_can;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_should;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_oprb_matches;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_oprb_can;
  wire  BufferedBroadcastAcquireTracker_3_1_io_alloc_oprb_should;
  wire  outer_arb_clk;
  wire  outer_arb_reset;
  wire  outer_arb_io_in_0_acquire_ready;
  wire  outer_arb_io_in_0_acquire_valid;
  wire [25:0] outer_arb_io_in_0_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_0_acquire_bits_addr_beat;
  wire  outer_arb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_0_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_0_acquire_bits_union;
  wire [63:0] outer_arb_io_in_0_acquire_bits_data;
  wire  outer_arb_io_in_0_probe_ready;
  wire  outer_arb_io_in_0_probe_valid;
  wire [25:0] outer_arb_io_in_0_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_0_probe_bits_p_type;
  wire  outer_arb_io_in_0_release_ready;
  wire  outer_arb_io_in_0_release_valid;
  wire [2:0] outer_arb_io_in_0_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_0_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_0_release_bits_client_xact_id;
  wire  outer_arb_io_in_0_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_0_release_bits_r_type;
  wire [63:0] outer_arb_io_in_0_release_bits_data;
  wire  outer_arb_io_in_0_grant_ready;
  wire  outer_arb_io_in_0_grant_valid;
  wire [2:0] outer_arb_io_in_0_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_0_grant_bits_client_xact_id;
  wire  outer_arb_io_in_0_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_0_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_0_grant_bits_data;
  wire  outer_arb_io_in_0_grant_bits_manager_id;
  wire  outer_arb_io_in_0_finish_ready;
  wire  outer_arb_io_in_0_finish_valid;
  wire  outer_arb_io_in_0_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_0_finish_bits_manager_id;
  wire  outer_arb_io_in_1_acquire_ready;
  wire  outer_arb_io_in_1_acquire_valid;
  wire [25:0] outer_arb_io_in_1_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_1_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_1_acquire_bits_addr_beat;
  wire  outer_arb_io_in_1_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_1_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_1_acquire_bits_union;
  wire [63:0] outer_arb_io_in_1_acquire_bits_data;
  wire  outer_arb_io_in_1_probe_ready;
  wire  outer_arb_io_in_1_probe_valid;
  wire [25:0] outer_arb_io_in_1_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_1_probe_bits_p_type;
  wire  outer_arb_io_in_1_release_ready;
  wire  outer_arb_io_in_1_release_valid;
  wire [2:0] outer_arb_io_in_1_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_1_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_1_release_bits_client_xact_id;
  wire  outer_arb_io_in_1_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_1_release_bits_r_type;
  wire [63:0] outer_arb_io_in_1_release_bits_data;
  wire  outer_arb_io_in_1_grant_ready;
  wire  outer_arb_io_in_1_grant_valid;
  wire [2:0] outer_arb_io_in_1_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_1_grant_bits_client_xact_id;
  wire  outer_arb_io_in_1_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_1_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_1_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_1_grant_bits_data;
  wire  outer_arb_io_in_1_grant_bits_manager_id;
  wire  outer_arb_io_in_1_finish_ready;
  wire  outer_arb_io_in_1_finish_valid;
  wire  outer_arb_io_in_1_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_1_finish_bits_manager_id;
  wire  outer_arb_io_in_2_acquire_ready;
  wire  outer_arb_io_in_2_acquire_valid;
  wire [25:0] outer_arb_io_in_2_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_2_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_2_acquire_bits_addr_beat;
  wire  outer_arb_io_in_2_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_2_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_2_acquire_bits_union;
  wire [63:0] outer_arb_io_in_2_acquire_bits_data;
  wire  outer_arb_io_in_2_probe_ready;
  wire  outer_arb_io_in_2_probe_valid;
  wire [25:0] outer_arb_io_in_2_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_2_probe_bits_p_type;
  wire  outer_arb_io_in_2_release_ready;
  wire  outer_arb_io_in_2_release_valid;
  wire [2:0] outer_arb_io_in_2_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_2_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_2_release_bits_client_xact_id;
  wire  outer_arb_io_in_2_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_2_release_bits_r_type;
  wire [63:0] outer_arb_io_in_2_release_bits_data;
  wire  outer_arb_io_in_2_grant_ready;
  wire  outer_arb_io_in_2_grant_valid;
  wire [2:0] outer_arb_io_in_2_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_2_grant_bits_client_xact_id;
  wire  outer_arb_io_in_2_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_2_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_2_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_2_grant_bits_data;
  wire  outer_arb_io_in_2_grant_bits_manager_id;
  wire  outer_arb_io_in_2_finish_ready;
  wire  outer_arb_io_in_2_finish_valid;
  wire  outer_arb_io_in_2_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_2_finish_bits_manager_id;
  wire  outer_arb_io_in_3_acquire_ready;
  wire  outer_arb_io_in_3_acquire_valid;
  wire [25:0] outer_arb_io_in_3_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_3_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_3_acquire_bits_addr_beat;
  wire  outer_arb_io_in_3_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_3_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_3_acquire_bits_union;
  wire [63:0] outer_arb_io_in_3_acquire_bits_data;
  wire  outer_arb_io_in_3_probe_ready;
  wire  outer_arb_io_in_3_probe_valid;
  wire [25:0] outer_arb_io_in_3_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_3_probe_bits_p_type;
  wire  outer_arb_io_in_3_release_ready;
  wire  outer_arb_io_in_3_release_valid;
  wire [2:0] outer_arb_io_in_3_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_3_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_3_release_bits_client_xact_id;
  wire  outer_arb_io_in_3_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_3_release_bits_r_type;
  wire [63:0] outer_arb_io_in_3_release_bits_data;
  wire  outer_arb_io_in_3_grant_ready;
  wire  outer_arb_io_in_3_grant_valid;
  wire [2:0] outer_arb_io_in_3_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_3_grant_bits_client_xact_id;
  wire  outer_arb_io_in_3_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_3_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_3_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_3_grant_bits_data;
  wire  outer_arb_io_in_3_grant_bits_manager_id;
  wire  outer_arb_io_in_3_finish_ready;
  wire  outer_arb_io_in_3_finish_valid;
  wire  outer_arb_io_in_3_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_3_finish_bits_manager_id;
  wire  outer_arb_io_in_4_acquire_ready;
  wire  outer_arb_io_in_4_acquire_valid;
  wire [25:0] outer_arb_io_in_4_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_4_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_4_acquire_bits_addr_beat;
  wire  outer_arb_io_in_4_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_4_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_4_acquire_bits_union;
  wire [63:0] outer_arb_io_in_4_acquire_bits_data;
  wire  outer_arb_io_in_4_probe_ready;
  wire  outer_arb_io_in_4_probe_valid;
  wire [25:0] outer_arb_io_in_4_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_4_probe_bits_p_type;
  wire  outer_arb_io_in_4_release_ready;
  wire  outer_arb_io_in_4_release_valid;
  wire [2:0] outer_arb_io_in_4_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_4_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_4_release_bits_client_xact_id;
  wire  outer_arb_io_in_4_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_4_release_bits_r_type;
  wire [63:0] outer_arb_io_in_4_release_bits_data;
  wire  outer_arb_io_in_4_grant_ready;
  wire  outer_arb_io_in_4_grant_valid;
  wire [2:0] outer_arb_io_in_4_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_4_grant_bits_client_xact_id;
  wire  outer_arb_io_in_4_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_4_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_4_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_4_grant_bits_data;
  wire  outer_arb_io_in_4_grant_bits_manager_id;
  wire  outer_arb_io_in_4_finish_ready;
  wire  outer_arb_io_in_4_finish_valid;
  wire  outer_arb_io_in_4_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_4_finish_bits_manager_id;
  wire  outer_arb_io_out_acquire_ready;
  wire  outer_arb_io_out_acquire_valid;
  wire [25:0] outer_arb_io_out_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_out_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_out_acquire_bits_addr_beat;
  wire  outer_arb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_out_acquire_bits_a_type;
  wire [11:0] outer_arb_io_out_acquire_bits_union;
  wire [63:0] outer_arb_io_out_acquire_bits_data;
  wire  outer_arb_io_out_probe_ready;
  wire  outer_arb_io_out_probe_valid;
  wire [25:0] outer_arb_io_out_probe_bits_addr_block;
  wire [1:0] outer_arb_io_out_probe_bits_p_type;
  wire  outer_arb_io_out_release_ready;
  wire  outer_arb_io_out_release_valid;
  wire [2:0] outer_arb_io_out_release_bits_addr_beat;
  wire [25:0] outer_arb_io_out_release_bits_addr_block;
  wire [2:0] outer_arb_io_out_release_bits_client_xact_id;
  wire  outer_arb_io_out_release_bits_voluntary;
  wire [2:0] outer_arb_io_out_release_bits_r_type;
  wire [63:0] outer_arb_io_out_release_bits_data;
  wire  outer_arb_io_out_grant_ready;
  wire  outer_arb_io_out_grant_valid;
  wire [2:0] outer_arb_io_out_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_out_grant_bits_client_xact_id;
  wire  outer_arb_io_out_grant_bits_manager_xact_id;
  wire  outer_arb_io_out_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_out_grant_bits_g_type;
  wire [63:0] outer_arb_io_out_grant_bits_data;
  wire  outer_arb_io_out_grant_bits_manager_id;
  wire  outer_arb_io_out_finish_ready;
  wire  outer_arb_io_out_finish_valid;
  wire  outer_arb_io_out_finish_bits_manager_xact_id;
  wire  outer_arb_io_out_finish_bits_manager_id;
  wire  T_1287;
  wire  T_1288;
  wire  irel_vs_iacq_conflict;
  wire  T_1290;
  wire  T_1296_0;
  wire  T_1296_1;
  wire  T_1296_2;
  wire  T_1296_3;
  wire  T_1296_4;
  wire [1:0] T_1298;
  wire [1:0] T_1299;
  wire [2:0] T_1300;
  wire [4:0] T_1301;
  wire  T_1307_0;
  wire  T_1307_1;
  wire  T_1307_2;
  wire  T_1307_3;
  wire  T_1307_4;
  wire [1:0] T_1309;
  wire [1:0] T_1310;
  wire [2:0] T_1311;
  wire [4:0] T_1312;
  wire  T_1313;
  wire  T_1314;
  wire  T_1315;
  wire  T_1316;
  wire  T_1317;
  wire [4:0] T_1325;
  wire [4:0] T_1326;
  wire [4:0] T_1327;
  wire [4:0] T_1328;
  wire [4:0] T_1329;
  wire  T_1335_0;
  wire  T_1335_1;
  wire  T_1335_2;
  wire  T_1335_3;
  wire  T_1335_4;
  wire [1:0] T_1337;
  wire [1:0] T_1338;
  wire [2:0] T_1339;
  wire [4:0] T_1340;
  wire [4:0] GEN_5;
  wire  T_1342;
  wire  T_1344;
  wire [4:0] T_1346;
  wire [4:0] T_1347;
  wire  T_1349;
  wire  T_1350;
  wire  T_1353;
  wire  T_1354;
  wire  T_1355;
  wire  T_1356;
  wire  T_1359;
  wire  T_1360;
  wire  T_1361;
  wire  T_1364;
  wire  T_1365;
  wire  T_1366;
  wire  T_1369;
  wire  T_1370;
  wire  T_1371;
  wire  T_1374;
  wire  T_1375;
  wire  T_1376;
  wire  T_1382_0;
  wire  T_1382_1;
  wire  T_1382_2;
  wire  T_1382_3;
  wire  T_1382_4;
  wire [1:0] T_1384;
  wire [1:0] T_1385;
  wire [2:0] T_1386;
  wire [4:0] T_1387;
  wire  T_1393_0;
  wire  T_1393_1;
  wire  T_1393_2;
  wire  T_1393_3;
  wire  T_1393_4;
  wire [1:0] T_1395;
  wire [1:0] T_1396;
  wire [2:0] T_1397;
  wire [4:0] T_1398;
  wire  T_1399;
  wire  T_1400;
  wire  T_1401;
  wire  T_1402;
  wire  T_1403;
  wire [4:0] T_1411;
  wire [4:0] T_1412;
  wire [4:0] T_1413;
  wire [4:0] T_1414;
  wire [4:0] T_1415;
  wire  T_1421_0;
  wire  T_1421_1;
  wire  T_1421_2;
  wire  T_1421_3;
  wire  T_1421_4;
  wire [1:0] T_1423;
  wire [1:0] T_1424;
  wire [2:0] T_1425;
  wire [4:0] T_1426;
  wire  T_1428;
  wire  T_1430;
  wire [4:0] T_1433;
  wire [4:0] T_1434;
  wire  T_1436;
  wire  T_1441;
  wire  T_1442;
  wire  T_1446;
  wire  T_1447;
  wire  T_1451;
  wire  T_1452;
  wire  T_1456;
  wire  T_1457;
  wire  T_1461;
  wire  T_1462;
  wire  LockingRRArbiter_7_1_clk;
  wire  LockingRRArbiter_7_1_reset;
  wire  LockingRRArbiter_7_1_io_in_0_ready;
  wire  LockingRRArbiter_7_1_io_in_0_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_0_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_0_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_0_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_1_ready;
  wire  LockingRRArbiter_7_1_io_in_1_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_1_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_1_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_1_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_2_ready;
  wire  LockingRRArbiter_7_1_io_in_2_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_2_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_2_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_2_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_3_ready;
  wire  LockingRRArbiter_7_1_io_in_3_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_3_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_3_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_3_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_4_ready;
  wire  LockingRRArbiter_7_1_io_in_4_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_4_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_4_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_4_bits_client_id;
  wire  LockingRRArbiter_7_1_io_out_ready;
  wire  LockingRRArbiter_7_1_io_out_valid;
  wire [25:0] LockingRRArbiter_7_1_io_out_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_out_bits_p_type;
  wire  LockingRRArbiter_7_1_io_out_bits_client_id;
  wire [2:0] LockingRRArbiter_7_1_io_chosen;
  wire  LockingRRArbiter_8_1_clk;
  wire  LockingRRArbiter_8_1_reset;
  wire  LockingRRArbiter_8_1_io_in_0_ready;
  wire  LockingRRArbiter_8_1_io_in_0_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_0_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_0_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_0_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_0_bits_data;
  wire  LockingRRArbiter_8_1_io_in_0_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_1_ready;
  wire  LockingRRArbiter_8_1_io_in_1_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_1_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_1_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_1_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_1_bits_data;
  wire  LockingRRArbiter_8_1_io_in_1_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_2_ready;
  wire  LockingRRArbiter_8_1_io_in_2_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_2_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_2_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_2_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_2_bits_data;
  wire  LockingRRArbiter_8_1_io_in_2_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_3_ready;
  wire  LockingRRArbiter_8_1_io_in_3_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_3_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_3_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_3_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_3_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_3_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_3_bits_data;
  wire  LockingRRArbiter_8_1_io_in_3_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_4_ready;
  wire  LockingRRArbiter_8_1_io_in_4_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_4_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_4_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_4_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_4_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_4_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_4_bits_data;
  wire  LockingRRArbiter_8_1_io_in_4_bits_client_id;
  wire  LockingRRArbiter_8_1_io_out_ready;
  wire  LockingRRArbiter_8_1_io_out_valid;
  wire [2:0] LockingRRArbiter_8_1_io_out_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_out_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_out_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_out_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_out_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_out_bits_data;
  wire  LockingRRArbiter_8_1_io_out_bits_client_id;
  wire [2:0] LockingRRArbiter_8_1_io_chosen;
  wire [2:0] GEN_9;
  wire  T_1465;
  wire  T_1466;
  wire [2:0] GEN_10;
  wire  T_1468;
  wire  T_1469;
  wire [2:0] GEN_11;
  wire  T_1471;
  wire  T_1472;
  wire [2:0] GEN_12;
  wire  T_1474;
  wire  T_1475;
  wire  T_1477;
  wire  T_1478;
  wire  T_1484_0;
  wire  T_1484_1;
  wire  T_1484_2;
  wire  T_1484_3;
  wire  T_1484_4;
  wire  GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  reg  GEN_6;
  reg [31:0] GEN_15;
  reg  GEN_7;
  reg [31:0] GEN_16;
  reg  GEN_8;
  reg [31:0] GEN_17;
  reg  GEN_13;
  reg [31:0] GEN_18;
  reg  GEN_14;
  reg [31:0] GEN_19;
  BufferedBroadcastVoluntaryReleaseTracker BufferedBroadcastVoluntaryReleaseTracker_1 (
    .clk(BufferedBroadcastVoluntaryReleaseTracker_1_clk),
    .reset(BufferedBroadcastVoluntaryReleaseTracker_1_reset),
    .io_inner_acquire_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_ready),
    .io_inner_grant_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_ready),
    .io_inner_finish_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_ready),
    .io_inner_probe_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_ready),
    .io_inner_release_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_client_id),
    .io_incoherent_0(BufferedBroadcastVoluntaryReleaseTracker_1_io_incoherent_0),
    .io_outer_acquire_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_ready),
    .io_outer_probe_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_ready),
    .io_outer_release_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_data),
    .io_outer_grant_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_ready),
    .io_outer_grant_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_ready),
    .io_outer_finish_valid(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_matches),
    .io_alloc_iacq_can(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_can),
    .io_alloc_iacq_should(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_should),
    .io_alloc_irel_matches(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_matches),
    .io_alloc_irel_can(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_can),
    .io_alloc_irel_should(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_should),
    .io_alloc_oprb_matches(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_oprb_matches),
    .io_alloc_oprb_can(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_oprb_can),
    .io_alloc_oprb_should(BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_oprb_should)
  );
  BufferedBroadcastAcquireTracker BufferedBroadcastAcquireTracker_4 (
    .clk(BufferedBroadcastAcquireTracker_4_clk),
    .reset(BufferedBroadcastAcquireTracker_4_reset),
    .io_inner_acquire_ready(BufferedBroadcastAcquireTracker_4_io_inner_acquire_ready),
    .io_inner_acquire_valid(BufferedBroadcastAcquireTracker_4_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BufferedBroadcastAcquireTracker_4_io_inner_grant_ready),
    .io_inner_grant_valid(BufferedBroadcastAcquireTracker_4_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BufferedBroadcastAcquireTracker_4_io_inner_finish_ready),
    .io_inner_finish_valid(BufferedBroadcastAcquireTracker_4_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BufferedBroadcastAcquireTracker_4_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BufferedBroadcastAcquireTracker_4_io_inner_probe_ready),
    .io_inner_probe_valid(BufferedBroadcastAcquireTracker_4_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BufferedBroadcastAcquireTracker_4_io_inner_release_ready),
    .io_inner_release_valid(BufferedBroadcastAcquireTracker_4_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BufferedBroadcastAcquireTracker_4_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BufferedBroadcastAcquireTracker_4_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BufferedBroadcastAcquireTracker_4_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BufferedBroadcastAcquireTracker_4_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BufferedBroadcastAcquireTracker_4_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BufferedBroadcastAcquireTracker_4_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BufferedBroadcastAcquireTracker_4_io_inner_release_bits_client_id),
    .io_incoherent_0(BufferedBroadcastAcquireTracker_4_io_incoherent_0),
    .io_outer_acquire_ready(BufferedBroadcastAcquireTracker_4_io_outer_acquire_ready),
    .io_outer_acquire_valid(BufferedBroadcastAcquireTracker_4_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_data),
    .io_outer_probe_ready(BufferedBroadcastAcquireTracker_4_io_outer_probe_ready),
    .io_outer_probe_valid(BufferedBroadcastAcquireTracker_4_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(BufferedBroadcastAcquireTracker_4_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(BufferedBroadcastAcquireTracker_4_io_outer_probe_bits_p_type),
    .io_outer_release_ready(BufferedBroadcastAcquireTracker_4_io_outer_release_ready),
    .io_outer_release_valid(BufferedBroadcastAcquireTracker_4_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(BufferedBroadcastAcquireTracker_4_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(BufferedBroadcastAcquireTracker_4_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(BufferedBroadcastAcquireTracker_4_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(BufferedBroadcastAcquireTracker_4_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(BufferedBroadcastAcquireTracker_4_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(BufferedBroadcastAcquireTracker_4_io_outer_release_bits_data),
    .io_outer_grant_ready(BufferedBroadcastAcquireTracker_4_io_outer_grant_ready),
    .io_outer_grant_valid(BufferedBroadcastAcquireTracker_4_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(BufferedBroadcastAcquireTracker_4_io_outer_finish_ready),
    .io_outer_finish_valid(BufferedBroadcastAcquireTracker_4_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(BufferedBroadcastAcquireTracker_4_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(BufferedBroadcastAcquireTracker_4_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(BufferedBroadcastAcquireTracker_4_io_alloc_iacq_matches),
    .io_alloc_iacq_can(BufferedBroadcastAcquireTracker_4_io_alloc_iacq_can),
    .io_alloc_iacq_should(BufferedBroadcastAcquireTracker_4_io_alloc_iacq_should),
    .io_alloc_irel_matches(BufferedBroadcastAcquireTracker_4_io_alloc_irel_matches),
    .io_alloc_irel_can(BufferedBroadcastAcquireTracker_4_io_alloc_irel_can),
    .io_alloc_irel_should(BufferedBroadcastAcquireTracker_4_io_alloc_irel_should),
    .io_alloc_oprb_matches(BufferedBroadcastAcquireTracker_4_io_alloc_oprb_matches),
    .io_alloc_oprb_can(BufferedBroadcastAcquireTracker_4_io_alloc_oprb_can),
    .io_alloc_oprb_should(BufferedBroadcastAcquireTracker_4_io_alloc_oprb_should)
  );
  BufferedBroadcastAcquireTracker_1 BufferedBroadcastAcquireTracker_1_1 (
    .clk(BufferedBroadcastAcquireTracker_1_1_clk),
    .reset(BufferedBroadcastAcquireTracker_1_1_reset),
    .io_inner_acquire_ready(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_ready),
    .io_inner_grant_valid(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BufferedBroadcastAcquireTracker_1_1_io_inner_finish_ready),
    .io_inner_finish_valid(BufferedBroadcastAcquireTracker_1_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BufferedBroadcastAcquireTracker_1_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BufferedBroadcastAcquireTracker_1_1_io_inner_probe_ready),
    .io_inner_probe_valid(BufferedBroadcastAcquireTracker_1_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BufferedBroadcastAcquireTracker_1_1_io_inner_release_ready),
    .io_inner_release_valid(BufferedBroadcastAcquireTracker_1_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_client_id),
    .io_incoherent_0(BufferedBroadcastAcquireTracker_1_1_io_incoherent_0),
    .io_outer_acquire_ready(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(BufferedBroadcastAcquireTracker_1_1_io_outer_probe_ready),
    .io_outer_probe_valid(BufferedBroadcastAcquireTracker_1_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(BufferedBroadcastAcquireTracker_1_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(BufferedBroadcastAcquireTracker_1_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(BufferedBroadcastAcquireTracker_1_1_io_outer_release_ready),
    .io_outer_release_valid(BufferedBroadcastAcquireTracker_1_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_data),
    .io_outer_grant_ready(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_ready),
    .io_outer_grant_valid(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(BufferedBroadcastAcquireTracker_1_1_io_outer_finish_ready),
    .io_outer_finish_valid(BufferedBroadcastAcquireTracker_1_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(BufferedBroadcastAcquireTracker_1_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(BufferedBroadcastAcquireTracker_1_1_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_matches),
    .io_alloc_iacq_can(BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_can),
    .io_alloc_iacq_should(BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_should),
    .io_alloc_irel_matches(BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_matches),
    .io_alloc_irel_can(BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_can),
    .io_alloc_irel_should(BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_should),
    .io_alloc_oprb_matches(BufferedBroadcastAcquireTracker_1_1_io_alloc_oprb_matches),
    .io_alloc_oprb_can(BufferedBroadcastAcquireTracker_1_1_io_alloc_oprb_can),
    .io_alloc_oprb_should(BufferedBroadcastAcquireTracker_1_1_io_alloc_oprb_should)
  );
  BufferedBroadcastAcquireTracker_2 BufferedBroadcastAcquireTracker_2_1 (
    .clk(BufferedBroadcastAcquireTracker_2_1_clk),
    .reset(BufferedBroadcastAcquireTracker_2_1_reset),
    .io_inner_acquire_ready(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_ready),
    .io_inner_grant_valid(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BufferedBroadcastAcquireTracker_2_1_io_inner_finish_ready),
    .io_inner_finish_valid(BufferedBroadcastAcquireTracker_2_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BufferedBroadcastAcquireTracker_2_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BufferedBroadcastAcquireTracker_2_1_io_inner_probe_ready),
    .io_inner_probe_valid(BufferedBroadcastAcquireTracker_2_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BufferedBroadcastAcquireTracker_2_1_io_inner_release_ready),
    .io_inner_release_valid(BufferedBroadcastAcquireTracker_2_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_client_id),
    .io_incoherent_0(BufferedBroadcastAcquireTracker_2_1_io_incoherent_0),
    .io_outer_acquire_ready(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(BufferedBroadcastAcquireTracker_2_1_io_outer_probe_ready),
    .io_outer_probe_valid(BufferedBroadcastAcquireTracker_2_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(BufferedBroadcastAcquireTracker_2_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(BufferedBroadcastAcquireTracker_2_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(BufferedBroadcastAcquireTracker_2_1_io_outer_release_ready),
    .io_outer_release_valid(BufferedBroadcastAcquireTracker_2_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_data),
    .io_outer_grant_ready(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_ready),
    .io_outer_grant_valid(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(BufferedBroadcastAcquireTracker_2_1_io_outer_finish_ready),
    .io_outer_finish_valid(BufferedBroadcastAcquireTracker_2_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(BufferedBroadcastAcquireTracker_2_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(BufferedBroadcastAcquireTracker_2_1_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_matches),
    .io_alloc_iacq_can(BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_can),
    .io_alloc_iacq_should(BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_should),
    .io_alloc_irel_matches(BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_matches),
    .io_alloc_irel_can(BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_can),
    .io_alloc_irel_should(BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_should),
    .io_alloc_oprb_matches(BufferedBroadcastAcquireTracker_2_1_io_alloc_oprb_matches),
    .io_alloc_oprb_can(BufferedBroadcastAcquireTracker_2_1_io_alloc_oprb_can),
    .io_alloc_oprb_should(BufferedBroadcastAcquireTracker_2_1_io_alloc_oprb_should)
  );
  BufferedBroadcastAcquireTracker_3 BufferedBroadcastAcquireTracker_3_1 (
    .clk(BufferedBroadcastAcquireTracker_3_1_clk),
    .reset(BufferedBroadcastAcquireTracker_3_1_reset),
    .io_inner_acquire_ready(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_ready),
    .io_inner_grant_valid(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BufferedBroadcastAcquireTracker_3_1_io_inner_finish_ready),
    .io_inner_finish_valid(BufferedBroadcastAcquireTracker_3_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BufferedBroadcastAcquireTracker_3_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BufferedBroadcastAcquireTracker_3_1_io_inner_probe_ready),
    .io_inner_probe_valid(BufferedBroadcastAcquireTracker_3_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BufferedBroadcastAcquireTracker_3_1_io_inner_release_ready),
    .io_inner_release_valid(BufferedBroadcastAcquireTracker_3_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_client_id),
    .io_incoherent_0(BufferedBroadcastAcquireTracker_3_1_io_incoherent_0),
    .io_outer_acquire_ready(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(BufferedBroadcastAcquireTracker_3_1_io_outer_probe_ready),
    .io_outer_probe_valid(BufferedBroadcastAcquireTracker_3_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(BufferedBroadcastAcquireTracker_3_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(BufferedBroadcastAcquireTracker_3_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(BufferedBroadcastAcquireTracker_3_1_io_outer_release_ready),
    .io_outer_release_valid(BufferedBroadcastAcquireTracker_3_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_data),
    .io_outer_grant_ready(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_ready),
    .io_outer_grant_valid(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(BufferedBroadcastAcquireTracker_3_1_io_outer_finish_ready),
    .io_outer_finish_valid(BufferedBroadcastAcquireTracker_3_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(BufferedBroadcastAcquireTracker_3_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(BufferedBroadcastAcquireTracker_3_1_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_matches),
    .io_alloc_iacq_can(BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_can),
    .io_alloc_iacq_should(BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_should),
    .io_alloc_irel_matches(BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_matches),
    .io_alloc_irel_can(BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_can),
    .io_alloc_irel_should(BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_should),
    .io_alloc_oprb_matches(BufferedBroadcastAcquireTracker_3_1_io_alloc_oprb_matches),
    .io_alloc_oprb_can(BufferedBroadcastAcquireTracker_3_1_io_alloc_oprb_can),
    .io_alloc_oprb_should(BufferedBroadcastAcquireTracker_3_1_io_alloc_oprb_should)
  );
  ClientTileLinkIOArbiter outer_arb (
    .clk(outer_arb_clk),
    .reset(outer_arb_reset),
    .io_in_0_acquire_ready(outer_arb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(outer_arb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(outer_arb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(outer_arb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(outer_arb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(outer_arb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(outer_arb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(outer_arb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(outer_arb_io_in_0_acquire_bits_data),
    .io_in_0_probe_ready(outer_arb_io_in_0_probe_ready),
    .io_in_0_probe_valid(outer_arb_io_in_0_probe_valid),
    .io_in_0_probe_bits_addr_block(outer_arb_io_in_0_probe_bits_addr_block),
    .io_in_0_probe_bits_p_type(outer_arb_io_in_0_probe_bits_p_type),
    .io_in_0_release_ready(outer_arb_io_in_0_release_ready),
    .io_in_0_release_valid(outer_arb_io_in_0_release_valid),
    .io_in_0_release_bits_addr_beat(outer_arb_io_in_0_release_bits_addr_beat),
    .io_in_0_release_bits_addr_block(outer_arb_io_in_0_release_bits_addr_block),
    .io_in_0_release_bits_client_xact_id(outer_arb_io_in_0_release_bits_client_xact_id),
    .io_in_0_release_bits_voluntary(outer_arb_io_in_0_release_bits_voluntary),
    .io_in_0_release_bits_r_type(outer_arb_io_in_0_release_bits_r_type),
    .io_in_0_release_bits_data(outer_arb_io_in_0_release_bits_data),
    .io_in_0_grant_ready(outer_arb_io_in_0_grant_ready),
    .io_in_0_grant_valid(outer_arb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(outer_arb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(outer_arb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(outer_arb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(outer_arb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(outer_arb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(outer_arb_io_in_0_grant_bits_data),
    .io_in_0_grant_bits_manager_id(outer_arb_io_in_0_grant_bits_manager_id),
    .io_in_0_finish_ready(outer_arb_io_in_0_finish_ready),
    .io_in_0_finish_valid(outer_arb_io_in_0_finish_valid),
    .io_in_0_finish_bits_manager_xact_id(outer_arb_io_in_0_finish_bits_manager_xact_id),
    .io_in_0_finish_bits_manager_id(outer_arb_io_in_0_finish_bits_manager_id),
    .io_in_1_acquire_ready(outer_arb_io_in_1_acquire_ready),
    .io_in_1_acquire_valid(outer_arb_io_in_1_acquire_valid),
    .io_in_1_acquire_bits_addr_block(outer_arb_io_in_1_acquire_bits_addr_block),
    .io_in_1_acquire_bits_client_xact_id(outer_arb_io_in_1_acquire_bits_client_xact_id),
    .io_in_1_acquire_bits_addr_beat(outer_arb_io_in_1_acquire_bits_addr_beat),
    .io_in_1_acquire_bits_is_builtin_type(outer_arb_io_in_1_acquire_bits_is_builtin_type),
    .io_in_1_acquire_bits_a_type(outer_arb_io_in_1_acquire_bits_a_type),
    .io_in_1_acquire_bits_union(outer_arb_io_in_1_acquire_bits_union),
    .io_in_1_acquire_bits_data(outer_arb_io_in_1_acquire_bits_data),
    .io_in_1_probe_ready(outer_arb_io_in_1_probe_ready),
    .io_in_1_probe_valid(outer_arb_io_in_1_probe_valid),
    .io_in_1_probe_bits_addr_block(outer_arb_io_in_1_probe_bits_addr_block),
    .io_in_1_probe_bits_p_type(outer_arb_io_in_1_probe_bits_p_type),
    .io_in_1_release_ready(outer_arb_io_in_1_release_ready),
    .io_in_1_release_valid(outer_arb_io_in_1_release_valid),
    .io_in_1_release_bits_addr_beat(outer_arb_io_in_1_release_bits_addr_beat),
    .io_in_1_release_bits_addr_block(outer_arb_io_in_1_release_bits_addr_block),
    .io_in_1_release_bits_client_xact_id(outer_arb_io_in_1_release_bits_client_xact_id),
    .io_in_1_release_bits_voluntary(outer_arb_io_in_1_release_bits_voluntary),
    .io_in_1_release_bits_r_type(outer_arb_io_in_1_release_bits_r_type),
    .io_in_1_release_bits_data(outer_arb_io_in_1_release_bits_data),
    .io_in_1_grant_ready(outer_arb_io_in_1_grant_ready),
    .io_in_1_grant_valid(outer_arb_io_in_1_grant_valid),
    .io_in_1_grant_bits_addr_beat(outer_arb_io_in_1_grant_bits_addr_beat),
    .io_in_1_grant_bits_client_xact_id(outer_arb_io_in_1_grant_bits_client_xact_id),
    .io_in_1_grant_bits_manager_xact_id(outer_arb_io_in_1_grant_bits_manager_xact_id),
    .io_in_1_grant_bits_is_builtin_type(outer_arb_io_in_1_grant_bits_is_builtin_type),
    .io_in_1_grant_bits_g_type(outer_arb_io_in_1_grant_bits_g_type),
    .io_in_1_grant_bits_data(outer_arb_io_in_1_grant_bits_data),
    .io_in_1_grant_bits_manager_id(outer_arb_io_in_1_grant_bits_manager_id),
    .io_in_1_finish_ready(outer_arb_io_in_1_finish_ready),
    .io_in_1_finish_valid(outer_arb_io_in_1_finish_valid),
    .io_in_1_finish_bits_manager_xact_id(outer_arb_io_in_1_finish_bits_manager_xact_id),
    .io_in_1_finish_bits_manager_id(outer_arb_io_in_1_finish_bits_manager_id),
    .io_in_2_acquire_ready(outer_arb_io_in_2_acquire_ready),
    .io_in_2_acquire_valid(outer_arb_io_in_2_acquire_valid),
    .io_in_2_acquire_bits_addr_block(outer_arb_io_in_2_acquire_bits_addr_block),
    .io_in_2_acquire_bits_client_xact_id(outer_arb_io_in_2_acquire_bits_client_xact_id),
    .io_in_2_acquire_bits_addr_beat(outer_arb_io_in_2_acquire_bits_addr_beat),
    .io_in_2_acquire_bits_is_builtin_type(outer_arb_io_in_2_acquire_bits_is_builtin_type),
    .io_in_2_acquire_bits_a_type(outer_arb_io_in_2_acquire_bits_a_type),
    .io_in_2_acquire_bits_union(outer_arb_io_in_2_acquire_bits_union),
    .io_in_2_acquire_bits_data(outer_arb_io_in_2_acquire_bits_data),
    .io_in_2_probe_ready(outer_arb_io_in_2_probe_ready),
    .io_in_2_probe_valid(outer_arb_io_in_2_probe_valid),
    .io_in_2_probe_bits_addr_block(outer_arb_io_in_2_probe_bits_addr_block),
    .io_in_2_probe_bits_p_type(outer_arb_io_in_2_probe_bits_p_type),
    .io_in_2_release_ready(outer_arb_io_in_2_release_ready),
    .io_in_2_release_valid(outer_arb_io_in_2_release_valid),
    .io_in_2_release_bits_addr_beat(outer_arb_io_in_2_release_bits_addr_beat),
    .io_in_2_release_bits_addr_block(outer_arb_io_in_2_release_bits_addr_block),
    .io_in_2_release_bits_client_xact_id(outer_arb_io_in_2_release_bits_client_xact_id),
    .io_in_2_release_bits_voluntary(outer_arb_io_in_2_release_bits_voluntary),
    .io_in_2_release_bits_r_type(outer_arb_io_in_2_release_bits_r_type),
    .io_in_2_release_bits_data(outer_arb_io_in_2_release_bits_data),
    .io_in_2_grant_ready(outer_arb_io_in_2_grant_ready),
    .io_in_2_grant_valid(outer_arb_io_in_2_grant_valid),
    .io_in_2_grant_bits_addr_beat(outer_arb_io_in_2_grant_bits_addr_beat),
    .io_in_2_grant_bits_client_xact_id(outer_arb_io_in_2_grant_bits_client_xact_id),
    .io_in_2_grant_bits_manager_xact_id(outer_arb_io_in_2_grant_bits_manager_xact_id),
    .io_in_2_grant_bits_is_builtin_type(outer_arb_io_in_2_grant_bits_is_builtin_type),
    .io_in_2_grant_bits_g_type(outer_arb_io_in_2_grant_bits_g_type),
    .io_in_2_grant_bits_data(outer_arb_io_in_2_grant_bits_data),
    .io_in_2_grant_bits_manager_id(outer_arb_io_in_2_grant_bits_manager_id),
    .io_in_2_finish_ready(outer_arb_io_in_2_finish_ready),
    .io_in_2_finish_valid(outer_arb_io_in_2_finish_valid),
    .io_in_2_finish_bits_manager_xact_id(outer_arb_io_in_2_finish_bits_manager_xact_id),
    .io_in_2_finish_bits_manager_id(outer_arb_io_in_2_finish_bits_manager_id),
    .io_in_3_acquire_ready(outer_arb_io_in_3_acquire_ready),
    .io_in_3_acquire_valid(outer_arb_io_in_3_acquire_valid),
    .io_in_3_acquire_bits_addr_block(outer_arb_io_in_3_acquire_bits_addr_block),
    .io_in_3_acquire_bits_client_xact_id(outer_arb_io_in_3_acquire_bits_client_xact_id),
    .io_in_3_acquire_bits_addr_beat(outer_arb_io_in_3_acquire_bits_addr_beat),
    .io_in_3_acquire_bits_is_builtin_type(outer_arb_io_in_3_acquire_bits_is_builtin_type),
    .io_in_3_acquire_bits_a_type(outer_arb_io_in_3_acquire_bits_a_type),
    .io_in_3_acquire_bits_union(outer_arb_io_in_3_acquire_bits_union),
    .io_in_3_acquire_bits_data(outer_arb_io_in_3_acquire_bits_data),
    .io_in_3_probe_ready(outer_arb_io_in_3_probe_ready),
    .io_in_3_probe_valid(outer_arb_io_in_3_probe_valid),
    .io_in_3_probe_bits_addr_block(outer_arb_io_in_3_probe_bits_addr_block),
    .io_in_3_probe_bits_p_type(outer_arb_io_in_3_probe_bits_p_type),
    .io_in_3_release_ready(outer_arb_io_in_3_release_ready),
    .io_in_3_release_valid(outer_arb_io_in_3_release_valid),
    .io_in_3_release_bits_addr_beat(outer_arb_io_in_3_release_bits_addr_beat),
    .io_in_3_release_bits_addr_block(outer_arb_io_in_3_release_bits_addr_block),
    .io_in_3_release_bits_client_xact_id(outer_arb_io_in_3_release_bits_client_xact_id),
    .io_in_3_release_bits_voluntary(outer_arb_io_in_3_release_bits_voluntary),
    .io_in_3_release_bits_r_type(outer_arb_io_in_3_release_bits_r_type),
    .io_in_3_release_bits_data(outer_arb_io_in_3_release_bits_data),
    .io_in_3_grant_ready(outer_arb_io_in_3_grant_ready),
    .io_in_3_grant_valid(outer_arb_io_in_3_grant_valid),
    .io_in_3_grant_bits_addr_beat(outer_arb_io_in_3_grant_bits_addr_beat),
    .io_in_3_grant_bits_client_xact_id(outer_arb_io_in_3_grant_bits_client_xact_id),
    .io_in_3_grant_bits_manager_xact_id(outer_arb_io_in_3_grant_bits_manager_xact_id),
    .io_in_3_grant_bits_is_builtin_type(outer_arb_io_in_3_grant_bits_is_builtin_type),
    .io_in_3_grant_bits_g_type(outer_arb_io_in_3_grant_bits_g_type),
    .io_in_3_grant_bits_data(outer_arb_io_in_3_grant_bits_data),
    .io_in_3_grant_bits_manager_id(outer_arb_io_in_3_grant_bits_manager_id),
    .io_in_3_finish_ready(outer_arb_io_in_3_finish_ready),
    .io_in_3_finish_valid(outer_arb_io_in_3_finish_valid),
    .io_in_3_finish_bits_manager_xact_id(outer_arb_io_in_3_finish_bits_manager_xact_id),
    .io_in_3_finish_bits_manager_id(outer_arb_io_in_3_finish_bits_manager_id),
    .io_in_4_acquire_ready(outer_arb_io_in_4_acquire_ready),
    .io_in_4_acquire_valid(outer_arb_io_in_4_acquire_valid),
    .io_in_4_acquire_bits_addr_block(outer_arb_io_in_4_acquire_bits_addr_block),
    .io_in_4_acquire_bits_client_xact_id(outer_arb_io_in_4_acquire_bits_client_xact_id),
    .io_in_4_acquire_bits_addr_beat(outer_arb_io_in_4_acquire_bits_addr_beat),
    .io_in_4_acquire_bits_is_builtin_type(outer_arb_io_in_4_acquire_bits_is_builtin_type),
    .io_in_4_acquire_bits_a_type(outer_arb_io_in_4_acquire_bits_a_type),
    .io_in_4_acquire_bits_union(outer_arb_io_in_4_acquire_bits_union),
    .io_in_4_acquire_bits_data(outer_arb_io_in_4_acquire_bits_data),
    .io_in_4_probe_ready(outer_arb_io_in_4_probe_ready),
    .io_in_4_probe_valid(outer_arb_io_in_4_probe_valid),
    .io_in_4_probe_bits_addr_block(outer_arb_io_in_4_probe_bits_addr_block),
    .io_in_4_probe_bits_p_type(outer_arb_io_in_4_probe_bits_p_type),
    .io_in_4_release_ready(outer_arb_io_in_4_release_ready),
    .io_in_4_release_valid(outer_arb_io_in_4_release_valid),
    .io_in_4_release_bits_addr_beat(outer_arb_io_in_4_release_bits_addr_beat),
    .io_in_4_release_bits_addr_block(outer_arb_io_in_4_release_bits_addr_block),
    .io_in_4_release_bits_client_xact_id(outer_arb_io_in_4_release_bits_client_xact_id),
    .io_in_4_release_bits_voluntary(outer_arb_io_in_4_release_bits_voluntary),
    .io_in_4_release_bits_r_type(outer_arb_io_in_4_release_bits_r_type),
    .io_in_4_release_bits_data(outer_arb_io_in_4_release_bits_data),
    .io_in_4_grant_ready(outer_arb_io_in_4_grant_ready),
    .io_in_4_grant_valid(outer_arb_io_in_4_grant_valid),
    .io_in_4_grant_bits_addr_beat(outer_arb_io_in_4_grant_bits_addr_beat),
    .io_in_4_grant_bits_client_xact_id(outer_arb_io_in_4_grant_bits_client_xact_id),
    .io_in_4_grant_bits_manager_xact_id(outer_arb_io_in_4_grant_bits_manager_xact_id),
    .io_in_4_grant_bits_is_builtin_type(outer_arb_io_in_4_grant_bits_is_builtin_type),
    .io_in_4_grant_bits_g_type(outer_arb_io_in_4_grant_bits_g_type),
    .io_in_4_grant_bits_data(outer_arb_io_in_4_grant_bits_data),
    .io_in_4_grant_bits_manager_id(outer_arb_io_in_4_grant_bits_manager_id),
    .io_in_4_finish_ready(outer_arb_io_in_4_finish_ready),
    .io_in_4_finish_valid(outer_arb_io_in_4_finish_valid),
    .io_in_4_finish_bits_manager_xact_id(outer_arb_io_in_4_finish_bits_manager_xact_id),
    .io_in_4_finish_bits_manager_id(outer_arb_io_in_4_finish_bits_manager_id),
    .io_out_acquire_ready(outer_arb_io_out_acquire_ready),
    .io_out_acquire_valid(outer_arb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(outer_arb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(outer_arb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(outer_arb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(outer_arb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(outer_arb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(outer_arb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(outer_arb_io_out_acquire_bits_data),
    .io_out_probe_ready(outer_arb_io_out_probe_ready),
    .io_out_probe_valid(outer_arb_io_out_probe_valid),
    .io_out_probe_bits_addr_block(outer_arb_io_out_probe_bits_addr_block),
    .io_out_probe_bits_p_type(outer_arb_io_out_probe_bits_p_type),
    .io_out_release_ready(outer_arb_io_out_release_ready),
    .io_out_release_valid(outer_arb_io_out_release_valid),
    .io_out_release_bits_addr_beat(outer_arb_io_out_release_bits_addr_beat),
    .io_out_release_bits_addr_block(outer_arb_io_out_release_bits_addr_block),
    .io_out_release_bits_client_xact_id(outer_arb_io_out_release_bits_client_xact_id),
    .io_out_release_bits_voluntary(outer_arb_io_out_release_bits_voluntary),
    .io_out_release_bits_r_type(outer_arb_io_out_release_bits_r_type),
    .io_out_release_bits_data(outer_arb_io_out_release_bits_data),
    .io_out_grant_ready(outer_arb_io_out_grant_ready),
    .io_out_grant_valid(outer_arb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(outer_arb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(outer_arb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(outer_arb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(outer_arb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(outer_arb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(outer_arb_io_out_grant_bits_data),
    .io_out_grant_bits_manager_id(outer_arb_io_out_grant_bits_manager_id),
    .io_out_finish_ready(outer_arb_io_out_finish_ready),
    .io_out_finish_valid(outer_arb_io_out_finish_valid),
    .io_out_finish_bits_manager_xact_id(outer_arb_io_out_finish_bits_manager_xact_id),
    .io_out_finish_bits_manager_id(outer_arb_io_out_finish_bits_manager_id)
  );
  LockingRRArbiter_7 LockingRRArbiter_7_1 (
    .clk(LockingRRArbiter_7_1_clk),
    .reset(LockingRRArbiter_7_1_reset),
    .io_in_0_ready(LockingRRArbiter_7_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_7_1_io_in_0_valid),
    .io_in_0_bits_addr_block(LockingRRArbiter_7_1_io_in_0_bits_addr_block),
    .io_in_0_bits_p_type(LockingRRArbiter_7_1_io_in_0_bits_p_type),
    .io_in_0_bits_client_id(LockingRRArbiter_7_1_io_in_0_bits_client_id),
    .io_in_1_ready(LockingRRArbiter_7_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_7_1_io_in_1_valid),
    .io_in_1_bits_addr_block(LockingRRArbiter_7_1_io_in_1_bits_addr_block),
    .io_in_1_bits_p_type(LockingRRArbiter_7_1_io_in_1_bits_p_type),
    .io_in_1_bits_client_id(LockingRRArbiter_7_1_io_in_1_bits_client_id),
    .io_in_2_ready(LockingRRArbiter_7_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_7_1_io_in_2_valid),
    .io_in_2_bits_addr_block(LockingRRArbiter_7_1_io_in_2_bits_addr_block),
    .io_in_2_bits_p_type(LockingRRArbiter_7_1_io_in_2_bits_p_type),
    .io_in_2_bits_client_id(LockingRRArbiter_7_1_io_in_2_bits_client_id),
    .io_in_3_ready(LockingRRArbiter_7_1_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_7_1_io_in_3_valid),
    .io_in_3_bits_addr_block(LockingRRArbiter_7_1_io_in_3_bits_addr_block),
    .io_in_3_bits_p_type(LockingRRArbiter_7_1_io_in_3_bits_p_type),
    .io_in_3_bits_client_id(LockingRRArbiter_7_1_io_in_3_bits_client_id),
    .io_in_4_ready(LockingRRArbiter_7_1_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_7_1_io_in_4_valid),
    .io_in_4_bits_addr_block(LockingRRArbiter_7_1_io_in_4_bits_addr_block),
    .io_in_4_bits_p_type(LockingRRArbiter_7_1_io_in_4_bits_p_type),
    .io_in_4_bits_client_id(LockingRRArbiter_7_1_io_in_4_bits_client_id),
    .io_out_ready(LockingRRArbiter_7_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_7_1_io_out_valid),
    .io_out_bits_addr_block(LockingRRArbiter_7_1_io_out_bits_addr_block),
    .io_out_bits_p_type(LockingRRArbiter_7_1_io_out_bits_p_type),
    .io_out_bits_client_id(LockingRRArbiter_7_1_io_out_bits_client_id),
    .io_chosen(LockingRRArbiter_7_1_io_chosen)
  );
  LockingRRArbiter_8 LockingRRArbiter_8_1 (
    .clk(LockingRRArbiter_8_1_clk),
    .reset(LockingRRArbiter_8_1_reset),
    .io_in_0_ready(LockingRRArbiter_8_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_8_1_io_in_0_valid),
    .io_in_0_bits_addr_beat(LockingRRArbiter_8_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_8_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(LockingRRArbiter_8_1_io_in_0_bits_g_type),
    .io_in_0_bits_data(LockingRRArbiter_8_1_io_in_0_bits_data),
    .io_in_0_bits_client_id(LockingRRArbiter_8_1_io_in_0_bits_client_id),
    .io_in_1_ready(LockingRRArbiter_8_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_8_1_io_in_1_valid),
    .io_in_1_bits_addr_beat(LockingRRArbiter_8_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_8_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(LockingRRArbiter_8_1_io_in_1_bits_g_type),
    .io_in_1_bits_data(LockingRRArbiter_8_1_io_in_1_bits_data),
    .io_in_1_bits_client_id(LockingRRArbiter_8_1_io_in_1_bits_client_id),
    .io_in_2_ready(LockingRRArbiter_8_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_8_1_io_in_2_valid),
    .io_in_2_bits_addr_beat(LockingRRArbiter_8_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_8_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(LockingRRArbiter_8_1_io_in_2_bits_g_type),
    .io_in_2_bits_data(LockingRRArbiter_8_1_io_in_2_bits_data),
    .io_in_2_bits_client_id(LockingRRArbiter_8_1_io_in_2_bits_client_id),
    .io_in_3_ready(LockingRRArbiter_8_1_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_8_1_io_in_3_valid),
    .io_in_3_bits_addr_beat(LockingRRArbiter_8_1_io_in_3_bits_addr_beat),
    .io_in_3_bits_client_xact_id(LockingRRArbiter_8_1_io_in_3_bits_client_xact_id),
    .io_in_3_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_3_bits_manager_xact_id),
    .io_in_3_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_g_type(LockingRRArbiter_8_1_io_in_3_bits_g_type),
    .io_in_3_bits_data(LockingRRArbiter_8_1_io_in_3_bits_data),
    .io_in_3_bits_client_id(LockingRRArbiter_8_1_io_in_3_bits_client_id),
    .io_in_4_ready(LockingRRArbiter_8_1_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_8_1_io_in_4_valid),
    .io_in_4_bits_addr_beat(LockingRRArbiter_8_1_io_in_4_bits_addr_beat),
    .io_in_4_bits_client_xact_id(LockingRRArbiter_8_1_io_in_4_bits_client_xact_id),
    .io_in_4_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_4_bits_manager_xact_id),
    .io_in_4_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_4_bits_is_builtin_type),
    .io_in_4_bits_g_type(LockingRRArbiter_8_1_io_in_4_bits_g_type),
    .io_in_4_bits_data(LockingRRArbiter_8_1_io_in_4_bits_data),
    .io_in_4_bits_client_id(LockingRRArbiter_8_1_io_in_4_bits_client_id),
    .io_out_ready(LockingRRArbiter_8_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_8_1_io_out_valid),
    .io_out_bits_addr_beat(LockingRRArbiter_8_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(LockingRRArbiter_8_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(LockingRRArbiter_8_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(LockingRRArbiter_8_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(LockingRRArbiter_8_1_io_out_bits_g_type),
    .io_out_bits_data(LockingRRArbiter_8_1_io_out_bits_data),
    .io_out_bits_client_id(LockingRRArbiter_8_1_io_out_bits_client_id),
    .io_chosen(LockingRRArbiter_8_1_io_chosen)
  );
  assign io_inner_acquire_ready = T_1350;
  assign io_inner_grant_valid = LockingRRArbiter_8_1_io_out_valid;
  assign io_inner_grant_bits_addr_beat = LockingRRArbiter_8_1_io_out_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = LockingRRArbiter_8_1_io_out_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = LockingRRArbiter_8_1_io_out_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = LockingRRArbiter_8_1_io_out_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = LockingRRArbiter_8_1_io_out_bits_g_type;
  assign io_inner_grant_bits_data = LockingRRArbiter_8_1_io_out_bits_data;
  assign io_inner_grant_bits_client_id = LockingRRArbiter_8_1_io_out_bits_client_id;
  assign io_inner_finish_ready = GEN_0;
  assign io_inner_probe_valid = LockingRRArbiter_7_1_io_out_valid;
  assign io_inner_probe_bits_addr_block = LockingRRArbiter_7_1_io_out_bits_addr_block;
  assign io_inner_probe_bits_p_type = LockingRRArbiter_7_1_io_out_bits_p_type;
  assign io_inner_probe_bits_client_id = LockingRRArbiter_7_1_io_out_bits_client_id;
  assign io_inner_release_ready = T_1436;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_outer_acquire_bits_addr_block = outer_arb_io_out_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_arb_io_out_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = outer_arb_io_out_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = outer_arb_io_out_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = outer_arb_io_out_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = outer_arb_io_out_acquire_bits_union;
  assign io_outer_acquire_bits_data = outer_arb_io_out_acquire_bits_data;
  assign io_outer_probe_ready = outer_arb_io_out_probe_ready;
  assign io_outer_release_valid = outer_arb_io_out_release_valid;
  assign io_outer_release_bits_addr_beat = outer_arb_io_out_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = outer_arb_io_out_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = outer_arb_io_out_release_bits_client_xact_id;
  assign io_outer_release_bits_voluntary = outer_arb_io_out_release_bits_voluntary;
  assign io_outer_release_bits_r_type = outer_arb_io_out_release_bits_r_type;
  assign io_outer_release_bits_data = outer_arb_io_out_release_bits_data;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_finish_valid = outer_arb_io_out_finish_valid;
  assign io_outer_finish_bits_manager_xact_id = outer_arb_io_out_finish_bits_manager_xact_id;
  assign io_outer_finish_bits_manager_id = outer_arb_io_out_finish_bits_manager_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_clk = clk;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_reset = reset;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_valid = T_1353;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_0_ready;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_valid = T_1466;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_0_ready;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_valid = io_inner_release_valid;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_data = io_inner_release_bits_data;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_incoherent_0 = io_incoherent_0;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_ready = outer_arb_io_in_0_acquire_ready;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_valid = outer_arb_io_in_0_probe_valid;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_bits_addr_block = outer_arb_io_in_0_probe_bits_addr_block;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_bits_p_type = outer_arb_io_in_0_probe_bits_p_type;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_ready = outer_arb_io_in_0_release_ready;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_valid = outer_arb_io_in_0_grant_valid;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_addr_beat = outer_arb_io_in_0_grant_bits_addr_beat;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_client_xact_id = outer_arb_io_in_0_grant_bits_client_xact_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_0_grant_bits_manager_xact_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_0_grant_bits_is_builtin_type;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_g_type = outer_arb_io_in_0_grant_bits_g_type;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_data = outer_arb_io_in_0_grant_bits_data;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_bits_manager_id = outer_arb_io_in_0_grant_bits_manager_id;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_ready = outer_arb_io_in_0_finish_ready;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_should = T_1356;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_should = T_1442;
  assign BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_oprb_should = GEN_6;
  assign BufferedBroadcastAcquireTracker_4_clk = clk;
  assign BufferedBroadcastAcquireTracker_4_reset = reset;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_valid = T_1353;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign BufferedBroadcastAcquireTracker_4_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BufferedBroadcastAcquireTracker_4_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_1_ready;
  assign BufferedBroadcastAcquireTracker_4_io_inner_finish_valid = T_1469;
  assign BufferedBroadcastAcquireTracker_4_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BufferedBroadcastAcquireTracker_4_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_1_ready;
  assign BufferedBroadcastAcquireTracker_4_io_inner_release_valid = io_inner_release_valid;
  assign BufferedBroadcastAcquireTracker_4_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_4_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_4_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_4_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BufferedBroadcastAcquireTracker_4_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BufferedBroadcastAcquireTracker_4_io_inner_release_bits_data = io_inner_release_bits_data;
  assign BufferedBroadcastAcquireTracker_4_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BufferedBroadcastAcquireTracker_4_io_incoherent_0 = io_incoherent_0;
  assign BufferedBroadcastAcquireTracker_4_io_outer_acquire_ready = outer_arb_io_in_1_acquire_ready;
  assign BufferedBroadcastAcquireTracker_4_io_outer_probe_valid = outer_arb_io_in_1_probe_valid;
  assign BufferedBroadcastAcquireTracker_4_io_outer_probe_bits_addr_block = outer_arb_io_in_1_probe_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_4_io_outer_probe_bits_p_type = outer_arb_io_in_1_probe_bits_p_type;
  assign BufferedBroadcastAcquireTracker_4_io_outer_release_ready = outer_arb_io_in_1_release_ready;
  assign BufferedBroadcastAcquireTracker_4_io_outer_grant_valid = outer_arb_io_in_1_grant_valid;
  assign BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_addr_beat = outer_arb_io_in_1_grant_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_client_xact_id = outer_arb_io_in_1_grant_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_1_grant_bits_manager_xact_id;
  assign BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_1_grant_bits_is_builtin_type;
  assign BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_g_type = outer_arb_io_in_1_grant_bits_g_type;
  assign BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_data = outer_arb_io_in_1_grant_bits_data;
  assign BufferedBroadcastAcquireTracker_4_io_outer_grant_bits_manager_id = outer_arb_io_in_1_grant_bits_manager_id;
  assign BufferedBroadcastAcquireTracker_4_io_outer_finish_ready = outer_arb_io_in_1_finish_ready;
  assign BufferedBroadcastAcquireTracker_4_io_alloc_iacq_should = T_1361;
  assign BufferedBroadcastAcquireTracker_4_io_alloc_irel_should = T_1447;
  assign BufferedBroadcastAcquireTracker_4_io_alloc_oprb_should = GEN_7;
  assign BufferedBroadcastAcquireTracker_1_1_clk = clk;
  assign BufferedBroadcastAcquireTracker_1_1_reset = reset;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_valid = T_1353;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_2_ready;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_finish_valid = T_1472;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_2_ready;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_release_valid = io_inner_release_valid;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_data = io_inner_release_bits_data;
  assign BufferedBroadcastAcquireTracker_1_1_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BufferedBroadcastAcquireTracker_1_1_io_incoherent_0 = io_incoherent_0;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_ready = outer_arb_io_in_2_acquire_ready;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_probe_valid = outer_arb_io_in_2_probe_valid;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_probe_bits_addr_block = outer_arb_io_in_2_probe_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_probe_bits_p_type = outer_arb_io_in_2_probe_bits_p_type;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_release_ready = outer_arb_io_in_2_release_ready;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_grant_valid = outer_arb_io_in_2_grant_valid;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_addr_beat = outer_arb_io_in_2_grant_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_client_xact_id = outer_arb_io_in_2_grant_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_2_grant_bits_manager_xact_id;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_2_grant_bits_is_builtin_type;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_g_type = outer_arb_io_in_2_grant_bits_g_type;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_data = outer_arb_io_in_2_grant_bits_data;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_grant_bits_manager_id = outer_arb_io_in_2_grant_bits_manager_id;
  assign BufferedBroadcastAcquireTracker_1_1_io_outer_finish_ready = outer_arb_io_in_2_finish_ready;
  assign BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_should = T_1366;
  assign BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_should = T_1452;
  assign BufferedBroadcastAcquireTracker_1_1_io_alloc_oprb_should = GEN_8;
  assign BufferedBroadcastAcquireTracker_2_1_clk = clk;
  assign BufferedBroadcastAcquireTracker_2_1_reset = reset;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_valid = T_1353;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_3_ready;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_finish_valid = T_1475;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_3_ready;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_release_valid = io_inner_release_valid;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_data = io_inner_release_bits_data;
  assign BufferedBroadcastAcquireTracker_2_1_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BufferedBroadcastAcquireTracker_2_1_io_incoherent_0 = io_incoherent_0;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_ready = outer_arb_io_in_3_acquire_ready;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_probe_valid = outer_arb_io_in_3_probe_valid;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_probe_bits_addr_block = outer_arb_io_in_3_probe_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_probe_bits_p_type = outer_arb_io_in_3_probe_bits_p_type;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_release_ready = outer_arb_io_in_3_release_ready;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_grant_valid = outer_arb_io_in_3_grant_valid;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_addr_beat = outer_arb_io_in_3_grant_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_client_xact_id = outer_arb_io_in_3_grant_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_3_grant_bits_manager_xact_id;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_3_grant_bits_is_builtin_type;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_g_type = outer_arb_io_in_3_grant_bits_g_type;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_data = outer_arb_io_in_3_grant_bits_data;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_grant_bits_manager_id = outer_arb_io_in_3_grant_bits_manager_id;
  assign BufferedBroadcastAcquireTracker_2_1_io_outer_finish_ready = outer_arb_io_in_3_finish_ready;
  assign BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_should = T_1371;
  assign BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_should = T_1457;
  assign BufferedBroadcastAcquireTracker_2_1_io_alloc_oprb_should = GEN_13;
  assign BufferedBroadcastAcquireTracker_3_1_clk = clk;
  assign BufferedBroadcastAcquireTracker_3_1_reset = reset;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_valid = T_1353;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_4_ready;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_finish_valid = T_1478;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_4_ready;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_release_valid = io_inner_release_valid;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_data = io_inner_release_bits_data;
  assign BufferedBroadcastAcquireTracker_3_1_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BufferedBroadcastAcquireTracker_3_1_io_incoherent_0 = io_incoherent_0;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_ready = outer_arb_io_in_4_acquire_ready;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_probe_valid = outer_arb_io_in_4_probe_valid;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_probe_bits_addr_block = outer_arb_io_in_4_probe_bits_addr_block;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_probe_bits_p_type = outer_arb_io_in_4_probe_bits_p_type;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_release_ready = outer_arb_io_in_4_release_ready;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_grant_valid = outer_arb_io_in_4_grant_valid;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_addr_beat = outer_arb_io_in_4_grant_bits_addr_beat;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_client_xact_id = outer_arb_io_in_4_grant_bits_client_xact_id;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_4_grant_bits_manager_xact_id;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_4_grant_bits_is_builtin_type;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_g_type = outer_arb_io_in_4_grant_bits_g_type;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_data = outer_arb_io_in_4_grant_bits_data;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_grant_bits_manager_id = outer_arb_io_in_4_grant_bits_manager_id;
  assign BufferedBroadcastAcquireTracker_3_1_io_outer_finish_ready = outer_arb_io_in_4_finish_ready;
  assign BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_should = T_1376;
  assign BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_should = T_1462;
  assign BufferedBroadcastAcquireTracker_3_1_io_alloc_oprb_should = GEN_14;
  assign outer_arb_clk = clk;
  assign outer_arb_reset = reset;
  assign outer_arb_io_in_0_acquire_valid = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_valid;
  assign outer_arb_io_in_0_acquire_bits_addr_block = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_0_acquire_bits_client_xact_id = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_0_acquire_bits_addr_beat = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_0_acquire_bits_is_builtin_type = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_0_acquire_bits_a_type = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_0_acquire_bits_union = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_union;
  assign outer_arb_io_in_0_acquire_bits_data = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_acquire_bits_data;
  assign outer_arb_io_in_0_probe_ready = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_probe_ready;
  assign outer_arb_io_in_0_release_valid = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_valid;
  assign outer_arb_io_in_0_release_bits_addr_beat = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_0_release_bits_addr_block = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_0_release_bits_client_xact_id = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_0_release_bits_voluntary = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_0_release_bits_r_type = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_r_type;
  assign outer_arb_io_in_0_release_bits_data = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_release_bits_data;
  assign outer_arb_io_in_0_grant_ready = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_grant_ready;
  assign outer_arb_io_in_0_finish_valid = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_valid;
  assign outer_arb_io_in_0_finish_bits_manager_xact_id = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_0_finish_bits_manager_id = BufferedBroadcastVoluntaryReleaseTracker_1_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_1_acquire_valid = BufferedBroadcastAcquireTracker_4_io_outer_acquire_valid;
  assign outer_arb_io_in_1_acquire_bits_addr_block = BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_1_acquire_bits_client_xact_id = BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_1_acquire_bits_addr_beat = BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_1_acquire_bits_is_builtin_type = BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_1_acquire_bits_a_type = BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_1_acquire_bits_union = BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_union;
  assign outer_arb_io_in_1_acquire_bits_data = BufferedBroadcastAcquireTracker_4_io_outer_acquire_bits_data;
  assign outer_arb_io_in_1_probe_ready = BufferedBroadcastAcquireTracker_4_io_outer_probe_ready;
  assign outer_arb_io_in_1_release_valid = BufferedBroadcastAcquireTracker_4_io_outer_release_valid;
  assign outer_arb_io_in_1_release_bits_addr_beat = BufferedBroadcastAcquireTracker_4_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_1_release_bits_addr_block = BufferedBroadcastAcquireTracker_4_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_1_release_bits_client_xact_id = BufferedBroadcastAcquireTracker_4_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_1_release_bits_voluntary = BufferedBroadcastAcquireTracker_4_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_1_release_bits_r_type = BufferedBroadcastAcquireTracker_4_io_outer_release_bits_r_type;
  assign outer_arb_io_in_1_release_bits_data = BufferedBroadcastAcquireTracker_4_io_outer_release_bits_data;
  assign outer_arb_io_in_1_grant_ready = BufferedBroadcastAcquireTracker_4_io_outer_grant_ready;
  assign outer_arb_io_in_1_finish_valid = BufferedBroadcastAcquireTracker_4_io_outer_finish_valid;
  assign outer_arb_io_in_1_finish_bits_manager_xact_id = BufferedBroadcastAcquireTracker_4_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_1_finish_bits_manager_id = BufferedBroadcastAcquireTracker_4_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_2_acquire_valid = BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_valid;
  assign outer_arb_io_in_2_acquire_bits_addr_block = BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_2_acquire_bits_client_xact_id = BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_2_acquire_bits_addr_beat = BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_2_acquire_bits_is_builtin_type = BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_2_acquire_bits_a_type = BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_2_acquire_bits_union = BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_union;
  assign outer_arb_io_in_2_acquire_bits_data = BufferedBroadcastAcquireTracker_1_1_io_outer_acquire_bits_data;
  assign outer_arb_io_in_2_probe_ready = BufferedBroadcastAcquireTracker_1_1_io_outer_probe_ready;
  assign outer_arb_io_in_2_release_valid = BufferedBroadcastAcquireTracker_1_1_io_outer_release_valid;
  assign outer_arb_io_in_2_release_bits_addr_beat = BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_2_release_bits_addr_block = BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_2_release_bits_client_xact_id = BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_2_release_bits_voluntary = BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_2_release_bits_r_type = BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_r_type;
  assign outer_arb_io_in_2_release_bits_data = BufferedBroadcastAcquireTracker_1_1_io_outer_release_bits_data;
  assign outer_arb_io_in_2_grant_ready = BufferedBroadcastAcquireTracker_1_1_io_outer_grant_ready;
  assign outer_arb_io_in_2_finish_valid = BufferedBroadcastAcquireTracker_1_1_io_outer_finish_valid;
  assign outer_arb_io_in_2_finish_bits_manager_xact_id = BufferedBroadcastAcquireTracker_1_1_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_2_finish_bits_manager_id = BufferedBroadcastAcquireTracker_1_1_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_3_acquire_valid = BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_valid;
  assign outer_arb_io_in_3_acquire_bits_addr_block = BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_3_acquire_bits_client_xact_id = BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_3_acquire_bits_addr_beat = BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_3_acquire_bits_is_builtin_type = BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_3_acquire_bits_a_type = BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_3_acquire_bits_union = BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_union;
  assign outer_arb_io_in_3_acquire_bits_data = BufferedBroadcastAcquireTracker_2_1_io_outer_acquire_bits_data;
  assign outer_arb_io_in_3_probe_ready = BufferedBroadcastAcquireTracker_2_1_io_outer_probe_ready;
  assign outer_arb_io_in_3_release_valid = BufferedBroadcastAcquireTracker_2_1_io_outer_release_valid;
  assign outer_arb_io_in_3_release_bits_addr_beat = BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_3_release_bits_addr_block = BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_3_release_bits_client_xact_id = BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_3_release_bits_voluntary = BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_3_release_bits_r_type = BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_r_type;
  assign outer_arb_io_in_3_release_bits_data = BufferedBroadcastAcquireTracker_2_1_io_outer_release_bits_data;
  assign outer_arb_io_in_3_grant_ready = BufferedBroadcastAcquireTracker_2_1_io_outer_grant_ready;
  assign outer_arb_io_in_3_finish_valid = BufferedBroadcastAcquireTracker_2_1_io_outer_finish_valid;
  assign outer_arb_io_in_3_finish_bits_manager_xact_id = BufferedBroadcastAcquireTracker_2_1_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_3_finish_bits_manager_id = BufferedBroadcastAcquireTracker_2_1_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_4_acquire_valid = BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_valid;
  assign outer_arb_io_in_4_acquire_bits_addr_block = BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_4_acquire_bits_client_xact_id = BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_4_acquire_bits_addr_beat = BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_4_acquire_bits_is_builtin_type = BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_4_acquire_bits_a_type = BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_4_acquire_bits_union = BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_union;
  assign outer_arb_io_in_4_acquire_bits_data = BufferedBroadcastAcquireTracker_3_1_io_outer_acquire_bits_data;
  assign outer_arb_io_in_4_probe_ready = BufferedBroadcastAcquireTracker_3_1_io_outer_probe_ready;
  assign outer_arb_io_in_4_release_valid = BufferedBroadcastAcquireTracker_3_1_io_outer_release_valid;
  assign outer_arb_io_in_4_release_bits_addr_beat = BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_4_release_bits_addr_block = BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_4_release_bits_client_xact_id = BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_4_release_bits_voluntary = BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_4_release_bits_r_type = BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_r_type;
  assign outer_arb_io_in_4_release_bits_data = BufferedBroadcastAcquireTracker_3_1_io_outer_release_bits_data;
  assign outer_arb_io_in_4_grant_ready = BufferedBroadcastAcquireTracker_3_1_io_outer_grant_ready;
  assign outer_arb_io_in_4_finish_valid = BufferedBroadcastAcquireTracker_3_1_io_outer_finish_valid;
  assign outer_arb_io_in_4_finish_bits_manager_xact_id = BufferedBroadcastAcquireTracker_3_1_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_4_finish_bits_manager_id = BufferedBroadcastAcquireTracker_3_1_io_outer_finish_bits_manager_id;
  assign outer_arb_io_out_acquire_ready = io_outer_acquire_ready;
  assign outer_arb_io_out_probe_valid = io_outer_probe_valid;
  assign outer_arb_io_out_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign outer_arb_io_out_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign outer_arb_io_out_release_ready = io_outer_release_ready;
  assign outer_arb_io_out_grant_valid = io_outer_grant_valid;
  assign outer_arb_io_out_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign outer_arb_io_out_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign outer_arb_io_out_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign outer_arb_io_out_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign outer_arb_io_out_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign outer_arb_io_out_grant_bits_data = io_outer_grant_bits_data;
  assign outer_arb_io_out_grant_bits_manager_id = io_outer_grant_bits_manager_id;
  assign outer_arb_io_out_finish_ready = io_outer_finish_ready;
  assign T_1287 = io_inner_acquire_valid & io_inner_release_valid;
  assign T_1288 = io_inner_release_bits_addr_block == io_inner_acquire_bits_addr_block;
  assign irel_vs_iacq_conflict = T_1287 & T_1288;
  assign T_1290 = irel_vs_iacq_conflict == 1'h0;
  assign T_1296_0 = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_acquire_ready;
  assign T_1296_1 = BufferedBroadcastAcquireTracker_4_io_inner_acquire_ready;
  assign T_1296_2 = BufferedBroadcastAcquireTracker_1_1_io_inner_acquire_ready;
  assign T_1296_3 = BufferedBroadcastAcquireTracker_2_1_io_inner_acquire_ready;
  assign T_1296_4 = BufferedBroadcastAcquireTracker_3_1_io_inner_acquire_ready;
  assign T_1298 = {T_1296_1,T_1296_0};
  assign T_1299 = {T_1296_4,T_1296_3};
  assign T_1300 = {T_1299,T_1296_2};
  assign T_1301 = {T_1300,T_1298};
  assign T_1307_0 = BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_can;
  assign T_1307_1 = BufferedBroadcastAcquireTracker_4_io_alloc_iacq_can;
  assign T_1307_2 = BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_can;
  assign T_1307_3 = BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_can;
  assign T_1307_4 = BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_can;
  assign T_1309 = {T_1307_1,T_1307_0};
  assign T_1310 = {T_1307_4,T_1307_3};
  assign T_1311 = {T_1310,T_1307_2};
  assign T_1312 = {T_1311,T_1309};
  assign T_1313 = T_1312[0];
  assign T_1314 = T_1312[1];
  assign T_1315 = T_1312[2];
  assign T_1316 = T_1312[3];
  assign T_1317 = T_1312[4];
  assign T_1325 = T_1317 ? 5'h10 : 5'h0;
  assign T_1326 = T_1316 ? 5'h8 : T_1325;
  assign T_1327 = T_1315 ? 5'h4 : T_1326;
  assign T_1328 = T_1314 ? 5'h2 : T_1327;
  assign T_1329 = T_1313 ? 5'h1 : T_1328;
  assign T_1335_0 = BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_iacq_matches;
  assign T_1335_1 = BufferedBroadcastAcquireTracker_4_io_alloc_iacq_matches;
  assign T_1335_2 = BufferedBroadcastAcquireTracker_1_1_io_alloc_iacq_matches;
  assign T_1335_3 = BufferedBroadcastAcquireTracker_2_1_io_alloc_iacq_matches;
  assign T_1335_4 = BufferedBroadcastAcquireTracker_3_1_io_alloc_iacq_matches;
  assign T_1337 = {T_1335_1,T_1335_0};
  assign T_1338 = {T_1335_4,T_1335_3};
  assign T_1339 = {T_1338,T_1335_2};
  assign T_1340 = {T_1339,T_1337};
  assign GEN_5 = {{4'd0}, 1'h0};
  assign T_1342 = T_1340 != GEN_5;
  assign T_1344 = T_1342 == 1'h0;
  assign T_1346 = T_1344 ? T_1312 : T_1340;
  assign T_1347 = T_1346 & T_1301;
  assign T_1349 = T_1347 != GEN_5;
  assign T_1350 = T_1349 & T_1290;
  assign T_1353 = io_inner_acquire_valid & T_1290;
  assign T_1354 = T_1329[0];
  assign T_1355 = T_1354 & T_1344;
  assign T_1356 = T_1355 & T_1290;
  assign T_1359 = T_1329[1];
  assign T_1360 = T_1359 & T_1344;
  assign T_1361 = T_1360 & T_1290;
  assign T_1364 = T_1329[2];
  assign T_1365 = T_1364 & T_1344;
  assign T_1366 = T_1365 & T_1290;
  assign T_1369 = T_1329[3];
  assign T_1370 = T_1369 & T_1344;
  assign T_1371 = T_1370 & T_1290;
  assign T_1374 = T_1329[4];
  assign T_1375 = T_1374 & T_1344;
  assign T_1376 = T_1375 & T_1290;
  assign T_1382_0 = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_release_ready;
  assign T_1382_1 = BufferedBroadcastAcquireTracker_4_io_inner_release_ready;
  assign T_1382_2 = BufferedBroadcastAcquireTracker_1_1_io_inner_release_ready;
  assign T_1382_3 = BufferedBroadcastAcquireTracker_2_1_io_inner_release_ready;
  assign T_1382_4 = BufferedBroadcastAcquireTracker_3_1_io_inner_release_ready;
  assign T_1384 = {T_1382_1,T_1382_0};
  assign T_1385 = {T_1382_4,T_1382_3};
  assign T_1386 = {T_1385,T_1382_2};
  assign T_1387 = {T_1386,T_1384};
  assign T_1393_0 = BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_can;
  assign T_1393_1 = BufferedBroadcastAcquireTracker_4_io_alloc_irel_can;
  assign T_1393_2 = BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_can;
  assign T_1393_3 = BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_can;
  assign T_1393_4 = BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_can;
  assign T_1395 = {T_1393_1,T_1393_0};
  assign T_1396 = {T_1393_4,T_1393_3};
  assign T_1397 = {T_1396,T_1393_2};
  assign T_1398 = {T_1397,T_1395};
  assign T_1399 = T_1398[0];
  assign T_1400 = T_1398[1];
  assign T_1401 = T_1398[2];
  assign T_1402 = T_1398[3];
  assign T_1403 = T_1398[4];
  assign T_1411 = T_1403 ? 5'h10 : 5'h0;
  assign T_1412 = T_1402 ? 5'h8 : T_1411;
  assign T_1413 = T_1401 ? 5'h4 : T_1412;
  assign T_1414 = T_1400 ? 5'h2 : T_1413;
  assign T_1415 = T_1399 ? 5'h1 : T_1414;
  assign T_1421_0 = BufferedBroadcastVoluntaryReleaseTracker_1_io_alloc_irel_matches;
  assign T_1421_1 = BufferedBroadcastAcquireTracker_4_io_alloc_irel_matches;
  assign T_1421_2 = BufferedBroadcastAcquireTracker_1_1_io_alloc_irel_matches;
  assign T_1421_3 = BufferedBroadcastAcquireTracker_2_1_io_alloc_irel_matches;
  assign T_1421_4 = BufferedBroadcastAcquireTracker_3_1_io_alloc_irel_matches;
  assign T_1423 = {T_1421_1,T_1421_0};
  assign T_1424 = {T_1421_4,T_1421_3};
  assign T_1425 = {T_1424,T_1421_2};
  assign T_1426 = {T_1425,T_1423};
  assign T_1428 = T_1426 != GEN_5;
  assign T_1430 = T_1428 == 1'h0;
  assign T_1433 = T_1430 ? T_1398 : T_1426;
  assign T_1434 = T_1433 & T_1387;
  assign T_1436 = T_1434 != GEN_5;
  assign T_1441 = T_1415[0];
  assign T_1442 = T_1441 & T_1430;
  assign T_1446 = T_1415[1];
  assign T_1447 = T_1446 & T_1430;
  assign T_1451 = T_1415[2];
  assign T_1452 = T_1451 & T_1430;
  assign T_1456 = T_1415[3];
  assign T_1457 = T_1456 & T_1430;
  assign T_1461 = T_1415[4];
  assign T_1462 = T_1461 & T_1430;
  assign LockingRRArbiter_7_1_clk = clk;
  assign LockingRRArbiter_7_1_reset = reset;
  assign LockingRRArbiter_7_1_io_in_0_valid = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_0_bits_addr_block = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_0_bits_p_type = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_0_bits_client_id = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_1_valid = BufferedBroadcastAcquireTracker_4_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_1_bits_addr_block = BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_1_bits_p_type = BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_1_bits_client_id = BufferedBroadcastAcquireTracker_4_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_2_valid = BufferedBroadcastAcquireTracker_1_1_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_2_bits_addr_block = BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_2_bits_p_type = BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_2_bits_client_id = BufferedBroadcastAcquireTracker_1_1_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_3_valid = BufferedBroadcastAcquireTracker_2_1_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_3_bits_addr_block = BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_3_bits_p_type = BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_3_bits_client_id = BufferedBroadcastAcquireTracker_2_1_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_4_valid = BufferedBroadcastAcquireTracker_3_1_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_4_bits_addr_block = BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_4_bits_p_type = BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_4_bits_client_id = BufferedBroadcastAcquireTracker_3_1_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_out_ready = io_inner_probe_ready;
  assign LockingRRArbiter_8_1_clk = clk;
  assign LockingRRArbiter_8_1_reset = reset;
  assign LockingRRArbiter_8_1_io_in_0_valid = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_0_bits_addr_beat = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_0_bits_client_xact_id = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_0_bits_g_type = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_0_bits_data = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_0_bits_client_id = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_1_valid = BufferedBroadcastAcquireTracker_4_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_1_bits_addr_beat = BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_1_bits_client_xact_id = BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id = BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type = BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_1_bits_g_type = BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_1_bits_data = BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_1_bits_client_id = BufferedBroadcastAcquireTracker_4_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_2_valid = BufferedBroadcastAcquireTracker_1_1_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_2_bits_addr_beat = BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_2_bits_client_xact_id = BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id = BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type = BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_2_bits_g_type = BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_2_bits_data = BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_2_bits_client_id = BufferedBroadcastAcquireTracker_1_1_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_3_valid = BufferedBroadcastAcquireTracker_2_1_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_3_bits_addr_beat = BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_3_bits_client_xact_id = BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_3_bits_manager_xact_id = BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_3_bits_is_builtin_type = BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_3_bits_g_type = BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_3_bits_data = BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_3_bits_client_id = BufferedBroadcastAcquireTracker_2_1_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_4_valid = BufferedBroadcastAcquireTracker_3_1_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_4_bits_addr_beat = BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_4_bits_client_xact_id = BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_4_bits_manager_xact_id = BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_4_bits_is_builtin_type = BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_4_bits_g_type = BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_4_bits_data = BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_4_bits_client_id = BufferedBroadcastAcquireTracker_3_1_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_out_ready = io_inner_grant_ready;
  assign GEN_9 = {{2'd0}, 1'h0};
  assign T_1465 = io_inner_finish_bits_manager_xact_id == GEN_9;
  assign T_1466 = io_inner_finish_valid & T_1465;
  assign GEN_10 = {{2'd0}, 1'h1};
  assign T_1468 = io_inner_finish_bits_manager_xact_id == GEN_10;
  assign T_1469 = io_inner_finish_valid & T_1468;
  assign GEN_11 = {{1'd0}, 2'h2};
  assign T_1471 = io_inner_finish_bits_manager_xact_id == GEN_11;
  assign T_1472 = io_inner_finish_valid & T_1471;
  assign GEN_12 = {{1'd0}, 2'h3};
  assign T_1474 = io_inner_finish_bits_manager_xact_id == GEN_12;
  assign T_1475 = io_inner_finish_valid & T_1474;
  assign T_1477 = io_inner_finish_bits_manager_xact_id == 3'h4;
  assign T_1478 = io_inner_finish_valid & T_1477;
  assign T_1484_0 = BufferedBroadcastVoluntaryReleaseTracker_1_io_inner_finish_ready;
  assign T_1484_1 = BufferedBroadcastAcquireTracker_4_io_inner_finish_ready;
  assign T_1484_2 = BufferedBroadcastAcquireTracker_1_1_io_inner_finish_ready;
  assign T_1484_3 = BufferedBroadcastAcquireTracker_2_1_io_inner_finish_ready;
  assign T_1484_4 = BufferedBroadcastAcquireTracker_3_1_io_inner_finish_ready;
  assign GEN_0 = GEN_4;
  assign GEN_1 = GEN_10 == io_inner_finish_bits_manager_xact_id ? T_1484_1 : T_1484_0;
  assign GEN_2 = GEN_11 == io_inner_finish_bits_manager_xact_id ? T_1484_2 : GEN_1;
  assign GEN_3 = GEN_12 == io_inner_finish_bits_manager_xact_id ? T_1484_3 : GEN_2;
  assign GEN_4 = 3'h4 == io_inner_finish_bits_manager_xact_id ? T_1484_4 : GEN_3;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  GEN_6 = GEN_15[0:0];
  GEN_16 = {1{$random}};
  GEN_7 = GEN_16[0:0];
  GEN_17 = {1{$random}};
  GEN_8 = GEN_17[0:0];
  GEN_18 = {1{$random}};
  GEN_13 = GEN_18[0:0];
  GEN_19 = {1{$random}};
  GEN_14 = GEN_19[0:0];
  end
`endif
endmodule
module MMIOTileLinkManager(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data
);
  wire  T_952;
  wire [2:0] T_961_0;
  wire  T_963;
  wire  T_966;
  wire  multibeat_fire;
  wire [2:0] GEN_43;
  wire  T_968;
  wire  multibeat_start;
  wire  T_970;
  wire  multibeat_end;
  reg [5:0] xact_pending;
  reg [31:0] GEN_54;
  wire [5:0] T_972;
  wire  T_973;
  wire  T_974;
  wire  T_975;
  wire  T_976;
  wire  T_977;
  wire [2:0] T_985;
  wire [2:0] T_986;
  wire [2:0] T_987;
  wire [2:0] T_988;
  wire [2:0] xact_id_sel;
  reg [2:0] xact_id_reg;
  reg [31:0] GEN_58;
  wire [2:0] GEN_4;
  reg  xact_multibeat;
  reg [31:0] GEN_59;
  wire [2:0] outer_xact_id;
  wire [5:0] GEN_44;
  wire  T_992;
  wire  xact_free;
  reg  xact_buffer_0_client_id;
  reg [31:0] GEN_60;
  reg [1:0] xact_buffer_0_client_xact_id;
  reg [31:0] GEN_61;
  reg  xact_buffer_1_client_id;
  reg [31:0] GEN_64;
  reg [1:0] xact_buffer_1_client_xact_id;
  reg [31:0] GEN_65;
  reg  xact_buffer_2_client_id;
  reg [31:0] GEN_66;
  reg [1:0] xact_buffer_2_client_xact_id;
  reg [31:0] GEN_67;
  reg  xact_buffer_3_client_id;
  reg [31:0] GEN_68;
  reg [1:0] xact_buffer_3_client_xact_id;
  reg [31:0] GEN_69;
  reg  xact_buffer_4_client_id;
  reg [31:0] GEN_70;
  reg [1:0] xact_buffer_4_client_xact_id;
  reg [31:0] GEN_71;
  reg  xact_buffer_5_client_id;
  reg [31:0] GEN_72;
  reg [1:0] xact_buffer_5_client_xact_id;
  reg [31:0] GEN_73;
  wire  T_1451;
  wire  T_1452;
  wire [2:0] T_1462_0;
  wire  T_1464;
  wire  T_1467;
  wire  T_1469;
  wire  T_1472;
  wire  T_1473;
  wire [3:0] GEN_45;
  wire [3:0] T_1475;
  wire [3:0] T_1477;
  wire [5:0] GEN_46;
  wire [5:0] T_1478;
  wire  T_1479;
  wire [7:0] GEN_47;
  wire [7:0] T_1481;
  wire [7:0] T_1483;
  wire [7:0] T_1484;
  wire [7:0] GEN_48;
  wire [7:0] T_1485;
  wire  T_1486;
  wire [2:0] T_1494_0;
  wire [3:0] GEN_49;
  wire  T_1496;
  wire [1:0] T_1504_0;
  wire [1:0] T_1504_1;
  wire [3:0] GEN_50;
  wire  T_1506;
  wire [3:0] GEN_51;
  wire  T_1507;
  wire  T_1510;
  wire  T_1511;
  wire  T_1514;
  wire  T_1516;
  wire  T_1517;
  wire  T_1518;
  wire [3:0] GEN_52;
  wire  T_1523;
  wire  T_1524;
  wire  T_1526;
  wire  T_1529;
  wire  T_1530;
  wire [7:0] T_1532;
  wire [7:0] T_1534;
  wire [7:0] T_1535;
  wire [7:0] T_1536;
  wire [2:0] T_1546_0;
  wire  T_1548;
  wire  T_1551;
  wire  T_1553;
  wire  T_1556;
  wire  T_1557;
  wire  GEN_0;
  wire  GEN_5;
  wire [2:0] GEN_55;
  wire  GEN_6;
  wire [2:0] GEN_56;
  wire  GEN_7;
  wire [2:0] GEN_57;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_1;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  wire [1:0] GEN_27;
  wire [1:0] GEN_28;
  wire [1:0] GEN_29;
  wire [1:0] GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_2;
  wire [1:0] GEN_62;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire [2:0] GEN_63;
  wire  GEN_36;
  wire  GEN_37;
  wire [1:0] GEN_3;
  wire [1:0] GEN_38;
  wire [1:0] GEN_39;
  wire [1:0] GEN_40;
  wire [1:0] GEN_41;
  wire [1:0] GEN_42;
  reg [25:0] GEN_17;
  reg [31:0] GEN_74;
  reg [1:0] GEN_24;
  reg [31:0] GEN_75;
  reg  GEN_53;
  reg [31:0] GEN_76;
  assign io_inner_acquire_ready = T_1451;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = GEN_3;
  assign io_inner_grant_bits_manager_xact_id = {{1'd0}, io_outer_grant_bits_client_xact_id};
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_client_id = GEN_2;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_17;
  assign io_inner_probe_bits_p_type = GEN_24;
  assign io_inner_probe_bits_client_id = GEN_53;
  assign io_inner_release_ready = 1'h0;
  assign io_outer_acquire_valid = T_1452;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_xact_id[1:0];
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign T_952 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_961_0 = 3'h3;
  assign T_963 = T_961_0 == io_outer_acquire_bits_a_type;
  assign T_966 = io_outer_acquire_bits_is_builtin_type & T_963;
  assign multibeat_fire = T_952 & T_966;
  assign GEN_43 = {{2'd0}, 1'h0};
  assign T_968 = io_outer_acquire_bits_addr_beat == GEN_43;
  assign multibeat_start = multibeat_fire & T_968;
  assign T_970 = io_outer_acquire_bits_addr_beat == 3'h7;
  assign multibeat_end = multibeat_fire & T_970;
  assign T_972 = ~ xact_pending;
  assign T_973 = T_972[0];
  assign T_974 = T_972[1];
  assign T_975 = T_972[2];
  assign T_976 = T_972[3];
  assign T_977 = T_972[4];
  assign T_985 = T_977 ? 3'h4 : 3'h5;
  assign T_986 = T_976 ? {{1'd0}, 2'h3} : T_985;
  assign T_987 = T_975 ? {{1'd0}, 2'h2} : T_986;
  assign T_988 = T_974 ? {{2'd0}, 1'h1} : T_987;
  assign xact_id_sel = T_973 ? {{2'd0}, 1'h0} : T_988;
  assign GEN_4 = multibeat_start ? xact_id_sel : xact_id_reg;
  assign outer_xact_id = xact_multibeat ? xact_id_reg : xact_id_sel;
  assign GEN_44 = {{5'd0}, 1'h0};
  assign T_992 = T_972 == GEN_44;
  assign xact_free = T_992 == 1'h0;
  assign T_1451 = io_outer_acquire_ready & xact_free;
  assign T_1452 = io_inner_acquire_valid & xact_free;
  assign T_1462_0 = 3'h3;
  assign T_1464 = T_1462_0 == io_outer_acquire_bits_a_type;
  assign T_1467 = io_outer_acquire_bits_is_builtin_type & T_1464;
  assign T_1469 = T_1467 == 1'h0;
  assign T_1472 = T_1469 | T_970;
  assign T_1473 = T_952 & T_1472;
  assign GEN_45 = {{3'd0}, 1'h1};
  assign T_1475 = GEN_45 << io_outer_acquire_bits_client_xact_id;
  assign T_1477 = T_1473 ? T_1475 : {{3'd0}, 1'h0};
  assign GEN_46 = {{2'd0}, T_1477};
  assign T_1478 = xact_pending | GEN_46;
  assign T_1479 = io_inner_finish_ready & io_inner_finish_valid;
  assign GEN_47 = {{7'd0}, 1'h1};
  assign T_1481 = GEN_47 << io_inner_finish_bits_manager_xact_id;
  assign T_1483 = T_1479 ? T_1481 : {{7'd0}, 1'h0};
  assign T_1484 = ~ T_1483;
  assign GEN_48 = {{2'd0}, T_1478};
  assign T_1485 = GEN_48 & T_1484;
  assign T_1486 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_1494_0 = 3'h5;
  assign GEN_49 = {{1'd0}, T_1494_0};
  assign T_1496 = GEN_49 == io_inner_grant_bits_g_type;
  assign T_1504_0 = 2'h0;
  assign T_1504_1 = 2'h1;
  assign GEN_50 = {{2'd0}, T_1504_0};
  assign T_1506 = GEN_50 == io_inner_grant_bits_g_type;
  assign GEN_51 = {{2'd0}, T_1504_1};
  assign T_1507 = GEN_51 == io_inner_grant_bits_g_type;
  assign T_1510 = T_1506 | T_1507;
  assign T_1511 = io_inner_grant_bits_is_builtin_type ? T_1496 : T_1510;
  assign T_1514 = T_1511 == 1'h0;
  assign T_1516 = io_inner_grant_bits_addr_beat == 3'h7;
  assign T_1517 = T_1514 | T_1516;
  assign T_1518 = T_1486 & T_1517;
  assign GEN_52 = {{1'd0}, 3'h0};
  assign T_1523 = io_inner_grant_bits_g_type == GEN_52;
  assign T_1524 = io_inner_grant_bits_is_builtin_type & T_1523;
  assign T_1526 = T_1524 == 1'h0;
  assign T_1529 = T_1526 == 1'h0;
  assign T_1530 = T_1518 & T_1529;
  assign T_1532 = GEN_47 << io_inner_grant_bits_manager_xact_id;
  assign T_1534 = T_1530 ? T_1532 : {{7'd0}, 1'h0};
  assign T_1535 = ~ T_1534;
  assign T_1536 = T_1485 & T_1535;
  assign T_1546_0 = 3'h3;
  assign T_1548 = T_1546_0 == io_outer_acquire_bits_a_type;
  assign T_1551 = io_outer_acquire_bits_is_builtin_type & T_1548;
  assign T_1553 = T_1551 == 1'h0;
  assign T_1556 = T_1553 | T_970;
  assign T_1557 = T_952 & T_1556;
  assign GEN_0 = io_inner_acquire_bits_client_id;
  assign GEN_5 = GEN_43 == outer_xact_id ? GEN_0 : xact_buffer_0_client_id;
  assign GEN_55 = {{2'd0}, 1'h1};
  assign GEN_6 = GEN_55 == outer_xact_id ? GEN_0 : xact_buffer_1_client_id;
  assign GEN_56 = {{1'd0}, 2'h2};
  assign GEN_7 = GEN_56 == outer_xact_id ? GEN_0 : xact_buffer_2_client_id;
  assign GEN_57 = {{1'd0}, 2'h3};
  assign GEN_8 = GEN_57 == outer_xact_id ? GEN_0 : xact_buffer_3_client_id;
  assign GEN_9 = 3'h4 == outer_xact_id ? GEN_0 : xact_buffer_4_client_id;
  assign GEN_10 = 3'h5 == outer_xact_id ? GEN_0 : xact_buffer_5_client_id;
  assign GEN_1 = io_inner_acquire_bits_client_xact_id;
  assign GEN_11 = GEN_43 == outer_xact_id ? GEN_1 : xact_buffer_0_client_xact_id;
  assign GEN_12 = GEN_55 == outer_xact_id ? GEN_1 : xact_buffer_1_client_xact_id;
  assign GEN_13 = GEN_56 == outer_xact_id ? GEN_1 : xact_buffer_2_client_xact_id;
  assign GEN_14 = GEN_57 == outer_xact_id ? GEN_1 : xact_buffer_3_client_xact_id;
  assign GEN_15 = 3'h4 == outer_xact_id ? GEN_1 : xact_buffer_4_client_xact_id;
  assign GEN_16 = 3'h5 == outer_xact_id ? GEN_1 : xact_buffer_5_client_xact_id;
  assign GEN_18 = T_1557 ? GEN_5 : xact_buffer_0_client_id;
  assign GEN_19 = T_1557 ? GEN_6 : xact_buffer_1_client_id;
  assign GEN_20 = T_1557 ? GEN_7 : xact_buffer_2_client_id;
  assign GEN_21 = T_1557 ? GEN_8 : xact_buffer_3_client_id;
  assign GEN_22 = T_1557 ? GEN_9 : xact_buffer_4_client_id;
  assign GEN_23 = T_1557 ? GEN_10 : xact_buffer_5_client_id;
  assign GEN_25 = T_1557 ? GEN_11 : xact_buffer_0_client_xact_id;
  assign GEN_26 = T_1557 ? GEN_12 : xact_buffer_1_client_xact_id;
  assign GEN_27 = T_1557 ? GEN_13 : xact_buffer_2_client_xact_id;
  assign GEN_28 = T_1557 ? GEN_14 : xact_buffer_3_client_xact_id;
  assign GEN_29 = T_1557 ? GEN_15 : xact_buffer_4_client_xact_id;
  assign GEN_30 = T_1557 ? GEN_16 : xact_buffer_5_client_xact_id;
  assign GEN_31 = multibeat_start ? 1'h1 : xact_multibeat;
  assign GEN_32 = multibeat_end ? 1'h0 : GEN_31;
  assign GEN_2 = GEN_37;
  assign GEN_62 = {{1'd0}, 1'h1};
  assign GEN_33 = GEN_62 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_id : xact_buffer_0_client_id;
  assign GEN_34 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_id : GEN_33;
  assign GEN_35 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_id : GEN_34;
  assign GEN_63 = {{1'd0}, io_outer_grant_bits_client_xact_id};
  assign GEN_36 = 3'h4 == GEN_63 ? xact_buffer_4_client_id : GEN_35;
  assign GEN_37 = 3'h5 == GEN_63 ? xact_buffer_5_client_id : GEN_36;
  assign GEN_3 = GEN_42;
  assign GEN_38 = GEN_62 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_xact_id : xact_buffer_0_client_xact_id;
  assign GEN_39 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_xact_id : GEN_38;
  assign GEN_40 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_xact_id : GEN_39;
  assign GEN_41 = 3'h4 == GEN_63 ? xact_buffer_4_client_xact_id : GEN_40;
  assign GEN_42 = 3'h5 == GEN_63 ? xact_buffer_5_client_xact_id : GEN_41;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_54 = {1{$random}};
  xact_pending = GEN_54[5:0];
  GEN_58 = {1{$random}};
  xact_id_reg = GEN_58[2:0];
  GEN_59 = {1{$random}};
  xact_multibeat = GEN_59[0:0];
  GEN_60 = {1{$random}};
  xact_buffer_0_client_id = GEN_60[0:0];
  GEN_61 = {1{$random}};
  xact_buffer_0_client_xact_id = GEN_61[1:0];
  GEN_64 = {1{$random}};
  xact_buffer_1_client_id = GEN_64[0:0];
  GEN_65 = {1{$random}};
  xact_buffer_1_client_xact_id = GEN_65[1:0];
  GEN_66 = {1{$random}};
  xact_buffer_2_client_id = GEN_66[0:0];
  GEN_67 = {1{$random}};
  xact_buffer_2_client_xact_id = GEN_67[1:0];
  GEN_68 = {1{$random}};
  xact_buffer_3_client_id = GEN_68[0:0];
  GEN_69 = {1{$random}};
  xact_buffer_3_client_xact_id = GEN_69[1:0];
  GEN_70 = {1{$random}};
  xact_buffer_4_client_id = GEN_70[0:0];
  GEN_71 = {1{$random}};
  xact_buffer_4_client_xact_id = GEN_71[1:0];
  GEN_72 = {1{$random}};
  xact_buffer_5_client_id = GEN_72[0:0];
  GEN_73 = {1{$random}};
  xact_buffer_5_client_xact_id = GEN_73[1:0];
  GEN_74 = {1{$random}};
  GEN_17 = GEN_74[25:0];
  GEN_75 = {1{$random}};
  GEN_24 = GEN_75[1:0];
  GEN_76 = {1{$random}};
  GEN_53 = GEN_76[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      xact_pending <= 6'h0;
    end else begin
      xact_pending <= T_1536[5:0];
    end
    if(1'h0) begin
    end else begin
      if(multibeat_start) begin
        if(T_973) begin
          xact_id_reg <= {{2'd0}, 1'h0};
        end else begin
          if(T_974) begin
            xact_id_reg <= {{2'd0}, 1'h1};
          end else begin
            if(T_975) begin
              xact_id_reg <= {{1'd0}, 2'h2};
            end else begin
              if(T_976) begin
                xact_id_reg <= {{1'd0}, 2'h3};
              end else begin
                if(T_977) begin
                  xact_id_reg <= 3'h4;
                end else begin
                  xact_id_reg <= 3'h5;
                end
              end
            end
          end
        end
      end
    end
    if(reset) begin
      xact_multibeat <= 1'h0;
    end else begin
      if(multibeat_end) begin
        xact_multibeat <= 1'h0;
      end else begin
        if(multibeat_start) begin
          xact_multibeat <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(GEN_43 == outer_xact_id) begin
          xact_buffer_0_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(GEN_43 == outer_xact_id) begin
          xact_buffer_0_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(GEN_55 == outer_xact_id) begin
          xact_buffer_1_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(GEN_55 == outer_xact_id) begin
          xact_buffer_1_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(GEN_56 == outer_xact_id) begin
          xact_buffer_2_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(GEN_56 == outer_xact_id) begin
          xact_buffer_2_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(GEN_57 == outer_xact_id) begin
          xact_buffer_3_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(GEN_57 == outer_xact_id) begin
          xact_buffer_3_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(3'h4 == outer_xact_id) begin
          xact_buffer_4_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(3'h4 == outer_xact_id) begin
          xact_buffer_4_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(3'h5 == outer_xact_id) begin
          xact_buffer_5_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1557) begin
        if(3'h5 == outer_xact_id) begin
          xact_buffer_5_client_xact_id <= GEN_1;
        end
      end
    end
  end
endmodule
module ClientUncachedTileLinkIOArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module TileLinkMemoryInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [2:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [2:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire  ClientUncachedTileLinkIOArbiter_1_1_clk;
  wire  ClientUncachedTileLinkIOArbiter_1_1_reset;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data;
  wire [25:0] T_3009;
  ClientUncachedTileLinkIOArbiter_1 ClientUncachedTileLinkIOArbiter_1_1 (
    .clk(ClientUncachedTileLinkIOArbiter_1_1_clk),
    .reset(ClientUncachedTileLinkIOArbiter_1_1_reset),
    .io_in_0_acquire_ready(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data),
    .io_out_acquire_ready(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready),
    .io_out_acquire_valid(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready),
    .io_out_grant_valid(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = T_3009;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_clk = clk;
  assign ClientUncachedTileLinkIOArbiter_1_1_reset = reset;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data = io_out_0_grant_bits_data;
  assign T_3009 = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block >> 1'h0;
endmodule
module LockingRRArbiter_9(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [2:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [11:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [2:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [11:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [2:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [11:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_8;
  wire [25:0] GEN_1;
  wire [25:0] GEN_9;
  wire [2:0] GEN_2;
  wire [2:0] GEN_10;
  wire [2:0] GEN_3;
  wire [2:0] GEN_11;
  wire  GEN_4;
  wire  GEN_12;
  wire [2:0] GEN_5;
  wire [2:0] GEN_13;
  wire [11:0] GEN_6;
  wire [11:0] GEN_14;
  wire [63:0] GEN_7;
  wire [63:0] GEN_15;
  reg [2:0] T_766;
  reg [31:0] GEN_24;
  reg  T_768;
  reg [31:0] GEN_25;
  wire [2:0] GEN_22;
  wire  T_770;
  wire [2:0] T_779_0;
  wire  T_781;
  wire  T_784;
  wire  T_785;
  wire  T_786;
  wire [2:0] GEN_23;
  wire [3:0] T_790;
  wire [2:0] T_791;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire  GEN_18;
  reg  lastGrant;
  reg [31:0] GEN_26;
  wire  GEN_19;
  wire  T_796;
  wire  T_798;
  wire  T_801;
  wire  T_805;
  wire  T_807;
  wire  T_811;
  wire  T_813;
  wire  T_814;
  wire  T_815;
  wire  T_818;
  wire  T_819;
  wire  GEN_20;
  wire  GEN_21;
  assign io_in_0_ready = T_815;
  assign io_in_1_ready = T_819;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_addr_beat = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_a_type = GEN_5;
  assign io_out_bits_union = GEN_6;
  assign io_out_bits_data = GEN_7;
  assign io_chosen = GEN_18;
  assign choice = GEN_21;
  assign GEN_0 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_2 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_3 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_4 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_5 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_6 = GEN_14;
  assign GEN_14 = io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_7 = GEN_15;
  assign GEN_15 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_22 = {{2'd0}, 1'h0};
  assign T_770 = T_766 != GEN_22;
  assign T_779_0 = 3'h3;
  assign T_781 = T_779_0 == io_out_bits_a_type;
  assign T_784 = io_out_bits_is_builtin_type & T_781;
  assign T_785 = io_out_ready & io_out_valid;
  assign T_786 = T_785 & T_784;
  assign GEN_23 = {{2'd0}, 1'h1};
  assign T_790 = T_766 + GEN_23;
  assign T_791 = T_790[2:0];
  assign GEN_16 = T_786 ? io_chosen : T_768;
  assign GEN_17 = T_786 ? T_791 : T_766;
  assign GEN_18 = T_770 ? T_768 : choice;
  assign GEN_19 = T_785 ? io_chosen : lastGrant;
  assign T_796 = 1'h1 > lastGrant;
  assign T_798 = io_in_1_valid & T_796;
  assign T_801 = T_798 | io_in_0_valid;
  assign T_805 = T_798 == 1'h0;
  assign T_807 = T_801 == 1'h0;
  assign T_811 = T_796 | T_807;
  assign T_813 = T_768 == 1'h0;
  assign T_814 = T_770 ? T_813 : T_805;
  assign T_815 = T_814 & io_out_ready;
  assign T_818 = T_770 ? T_768 : T_811;
  assign T_819 = T_818 & io_out_ready;
  assign GEN_20 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_21 = T_798 ? 1'h1 : GEN_20;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_24 = {1{$random}};
  T_766 = GEN_24[2:0];
  GEN_25 = {1{$random}};
  T_768 = GEN_25[0:0];
  GEN_26 = {1{$random}};
  lastGrant = GEN_26[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_766 <= 3'h0;
    end else begin
      if(T_786) begin
        T_766 <= T_791;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_786) begin
        T_768 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_785) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ReorderQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_data,
  input  [2:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [2:0] io_deq_tag,
  output  io_deq_data,
  output  io_deq_matches
);
  reg  roq_data [0:5];
  reg [31:0] GEN_15;
  wire  roq_data_T_104_data;
  wire [2:0] roq_data_T_104_addr;
  wire  roq_data_T_104_en;
  wire  roq_data_T_111_data;
  wire [2:0] roq_data_T_111_addr;
  wire  roq_data_T_111_mask;
  wire  roq_data_T_111_en;
  reg [2:0] roq_tags_0;
  reg [31:0] GEN_16;
  reg [2:0] roq_tags_1;
  reg [31:0] GEN_17;
  reg [2:0] roq_tags_2;
  reg [31:0] GEN_18;
  reg [2:0] roq_tags_3;
  reg [31:0] GEN_19;
  reg [2:0] roq_tags_4;
  reg [31:0] GEN_20;
  reg [2:0] roq_tags_5;
  reg [31:0] GEN_27;
  wire  T_50_0;
  wire  T_50_1;
  wire  T_50_2;
  wire  T_50_3;
  wire  T_50_4;
  wire  T_50_5;
  reg  roq_free_0;
  reg [31:0] GEN_40;
  reg  roq_free_1;
  reg [31:0] GEN_51;
  reg  roq_free_2;
  reg [31:0] GEN_52;
  reg  roq_free_3;
  reg [31:0] GEN_53;
  reg  roq_free_4;
  reg [31:0] GEN_54;
  reg  roq_free_5;
  reg [31:0] GEN_55;
  wire [2:0] T_61;
  wire [2:0] T_62;
  wire [2:0] T_63;
  wire [2:0] T_64;
  wire [2:0] roq_enq_addr;
  wire  T_65;
  wire  T_67;
  wire  T_68;
  wire  T_69;
  wire  T_71;
  wire  T_72;
  wire  T_73;
  wire  T_75;
  wire  T_76;
  wire  T_77;
  wire  T_79;
  wire  T_80;
  wire  T_81;
  wire  T_83;
  wire  T_84;
  wire  T_85;
  wire  T_87;
  wire  T_88;
  wire [2:0] T_95;
  wire [2:0] T_96;
  wire [2:0] T_97;
  wire [2:0] T_98;
  wire [2:0] roq_deq_addr;
  wire  T_99;
  wire  T_100;
  wire  T_101;
  wire  T_102;
  wire  T_103;
  wire  T_105;
  wire  T_106;
  wire  T_107;
  wire  T_108;
  wire  T_109;
  wire  T_110;
  wire [2:0] GEN_0;
  wire [2:0] GEN_47;
  wire [2:0] GEN_3;
  wire [2:0] GEN_48;
  wire [2:0] GEN_4;
  wire [2:0] GEN_49;
  wire [2:0] GEN_5;
  wire [2:0] GEN_50;
  wire [2:0] GEN_6;
  wire [2:0] GEN_7;
  wire [2:0] GEN_8;
  wire  GEN_1;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire [2:0] GEN_24;
  wire [2:0] GEN_25;
  wire [2:0] GEN_26;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_2;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  assign io_enq_ready = T_103;
  assign io_deq_data = roq_data_T_104_data;
  assign io_deq_matches = T_109;
  assign roq_data_T_104_addr = roq_deq_addr;
  assign roq_data_T_104_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_T_104_data = roq_data[roq_data_T_104_addr];
  `else
  assign roq_data_T_104_data = roq_data_T_104_addr >= 3'h6 ? $random : roq_data[roq_data_T_104_addr];
  `endif
  assign roq_data_T_111_data = io_enq_bits_data;
  assign roq_data_T_111_addr = roq_enq_addr;
  assign roq_data_T_111_mask = T_110;
  assign roq_data_T_111_en = T_110;
  assign T_50_0 = 1'h1;
  assign T_50_1 = 1'h1;
  assign T_50_2 = 1'h1;
  assign T_50_3 = 1'h1;
  assign T_50_4 = 1'h1;
  assign T_50_5 = 1'h1;
  assign T_61 = roq_free_4 ? 3'h4 : 3'h5;
  assign T_62 = roq_free_3 ? {{1'd0}, 2'h3} : T_61;
  assign T_63 = roq_free_2 ? {{1'd0}, 2'h2} : T_62;
  assign T_64 = roq_free_1 ? {{2'd0}, 1'h1} : T_63;
  assign roq_enq_addr = roq_free_0 ? {{2'd0}, 1'h0} : T_64;
  assign T_65 = roq_tags_0 == io_deq_tag;
  assign T_67 = roq_free_0 == 1'h0;
  assign T_68 = T_65 & T_67;
  assign T_69 = roq_tags_1 == io_deq_tag;
  assign T_71 = roq_free_1 == 1'h0;
  assign T_72 = T_69 & T_71;
  assign T_73 = roq_tags_2 == io_deq_tag;
  assign T_75 = roq_free_2 == 1'h0;
  assign T_76 = T_73 & T_75;
  assign T_77 = roq_tags_3 == io_deq_tag;
  assign T_79 = roq_free_3 == 1'h0;
  assign T_80 = T_77 & T_79;
  assign T_81 = roq_tags_4 == io_deq_tag;
  assign T_83 = roq_free_4 == 1'h0;
  assign T_84 = T_81 & T_83;
  assign T_85 = roq_tags_5 == io_deq_tag;
  assign T_87 = roq_free_5 == 1'h0;
  assign T_88 = T_85 & T_87;
  assign T_95 = T_84 ? 3'h4 : 3'h5;
  assign T_96 = T_80 ? {{1'd0}, 2'h3} : T_95;
  assign T_97 = T_76 ? {{1'd0}, 2'h2} : T_96;
  assign T_98 = T_72 ? {{2'd0}, 1'h1} : T_97;
  assign roq_deq_addr = T_68 ? {{2'd0}, 1'h0} : T_98;
  assign T_99 = roq_free_0 | roq_free_1;
  assign T_100 = T_99 | roq_free_2;
  assign T_101 = T_100 | roq_free_3;
  assign T_102 = T_101 | roq_free_4;
  assign T_103 = T_102 | roq_free_5;
  assign T_105 = T_68 | T_72;
  assign T_106 = T_105 | T_76;
  assign T_107 = T_106 | T_80;
  assign T_108 = T_107 | T_84;
  assign T_109 = T_108 | T_88;
  assign T_110 = io_enq_valid & io_enq_ready;
  assign GEN_0 = io_enq_bits_tag;
  assign GEN_47 = {{2'd0}, 1'h0};
  assign GEN_3 = GEN_47 == roq_enq_addr ? GEN_0 : roq_tags_0;
  assign GEN_48 = {{2'd0}, 1'h1};
  assign GEN_4 = GEN_48 == roq_enq_addr ? GEN_0 : roq_tags_1;
  assign GEN_49 = {{1'd0}, 2'h2};
  assign GEN_5 = GEN_49 == roq_enq_addr ? GEN_0 : roq_tags_2;
  assign GEN_50 = {{1'd0}, 2'h3};
  assign GEN_6 = GEN_50 == roq_enq_addr ? GEN_0 : roq_tags_3;
  assign GEN_7 = 3'h4 == roq_enq_addr ? GEN_0 : roq_tags_4;
  assign GEN_8 = 3'h5 == roq_enq_addr ? GEN_0 : roq_tags_5;
  assign GEN_1 = 1'h0;
  assign GEN_9 = GEN_47 == roq_enq_addr ? GEN_1 : roq_free_0;
  assign GEN_10 = GEN_48 == roq_enq_addr ? GEN_1 : roq_free_1;
  assign GEN_11 = GEN_49 == roq_enq_addr ? GEN_1 : roq_free_2;
  assign GEN_12 = GEN_50 == roq_enq_addr ? GEN_1 : roq_free_3;
  assign GEN_13 = 3'h4 == roq_enq_addr ? GEN_1 : roq_free_4;
  assign GEN_14 = 3'h5 == roq_enq_addr ? GEN_1 : roq_free_5;
  assign GEN_21 = T_110 ? GEN_3 : roq_tags_0;
  assign GEN_22 = T_110 ? GEN_4 : roq_tags_1;
  assign GEN_23 = T_110 ? GEN_5 : roq_tags_2;
  assign GEN_24 = T_110 ? GEN_6 : roq_tags_3;
  assign GEN_25 = T_110 ? GEN_7 : roq_tags_4;
  assign GEN_26 = T_110 ? GEN_8 : roq_tags_5;
  assign GEN_28 = T_110 ? GEN_9 : roq_free_0;
  assign GEN_29 = T_110 ? GEN_10 : roq_free_1;
  assign GEN_30 = T_110 ? GEN_11 : roq_free_2;
  assign GEN_31 = T_110 ? GEN_12 : roq_free_3;
  assign GEN_32 = T_110 ? GEN_13 : roq_free_4;
  assign GEN_33 = T_110 ? GEN_14 : roq_free_5;
  assign GEN_2 = 1'h1;
  assign GEN_34 = GEN_47 == roq_deq_addr ? GEN_2 : GEN_28;
  assign GEN_35 = GEN_48 == roq_deq_addr ? GEN_2 : GEN_29;
  assign GEN_36 = GEN_49 == roq_deq_addr ? GEN_2 : GEN_30;
  assign GEN_37 = GEN_50 == roq_deq_addr ? GEN_2 : GEN_31;
  assign GEN_38 = 3'h4 == roq_deq_addr ? GEN_2 : GEN_32;
  assign GEN_39 = 3'h5 == roq_deq_addr ? GEN_2 : GEN_33;
  assign GEN_41 = io_deq_valid ? GEN_34 : GEN_28;
  assign GEN_42 = io_deq_valid ? GEN_35 : GEN_29;
  assign GEN_43 = io_deq_valid ? GEN_36 : GEN_30;
  assign GEN_44 = io_deq_valid ? GEN_37 : GEN_31;
  assign GEN_45 = io_deq_valid ? GEN_38 : GEN_32;
  assign GEN_46 = io_deq_valid ? GEN_39 : GEN_33;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    roq_data[initvar] = GEN_15[0:0];
  GEN_16 = {1{$random}};
  roq_tags_0 = GEN_16[2:0];
  GEN_17 = {1{$random}};
  roq_tags_1 = GEN_17[2:0];
  GEN_18 = {1{$random}};
  roq_tags_2 = GEN_18[2:0];
  GEN_19 = {1{$random}};
  roq_tags_3 = GEN_19[2:0];
  GEN_20 = {1{$random}};
  roq_tags_4 = GEN_20[2:0];
  GEN_27 = {1{$random}};
  roq_tags_5 = GEN_27[2:0];
  GEN_40 = {1{$random}};
  roq_free_0 = GEN_40[0:0];
  GEN_51 = {1{$random}};
  roq_free_1 = GEN_51[0:0];
  GEN_52 = {1{$random}};
  roq_free_2 = GEN_52[0:0];
  GEN_53 = {1{$random}};
  roq_free_3 = GEN_53[0:0];
  GEN_54 = {1{$random}};
  roq_free_4 = GEN_54[0:0];
  GEN_55 = {1{$random}};
  roq_free_5 = GEN_55[0:0];
  end
`endif
  always @(posedge clk) begin
    if(roq_data_T_111_en & roq_data_T_111_mask) begin
      roq_data[roq_data_T_111_addr] <= roq_data_T_111_data;
    end
    if(1'h0) begin
    end else begin
      if(T_110) begin
        if(GEN_47 == roq_enq_addr) begin
          roq_tags_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_110) begin
        if(GEN_48 == roq_enq_addr) begin
          roq_tags_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_110) begin
        if(GEN_49 == roq_enq_addr) begin
          roq_tags_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_110) begin
        if(GEN_50 == roq_enq_addr) begin
          roq_tags_3 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_110) begin
        if(3'h4 == roq_enq_addr) begin
          roq_tags_4 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_110) begin
        if(3'h5 == roq_enq_addr) begin
          roq_tags_5 <= GEN_0;
        end
      end
    end
    if(reset) begin
      roq_free_0 <= T_50_0;
    end else begin
      if(io_deq_valid) begin
        if(GEN_47 == roq_deq_addr) begin
          roq_free_0 <= GEN_2;
        end else begin
          if(T_110) begin
            if(GEN_47 == roq_enq_addr) begin
              roq_free_0 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_110) begin
          if(GEN_47 == roq_enq_addr) begin
            roq_free_0 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_1 <= T_50_1;
    end else begin
      if(io_deq_valid) begin
        if(GEN_48 == roq_deq_addr) begin
          roq_free_1 <= GEN_2;
        end else begin
          if(T_110) begin
            if(GEN_48 == roq_enq_addr) begin
              roq_free_1 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_110) begin
          if(GEN_48 == roq_enq_addr) begin
            roq_free_1 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_2 <= T_50_2;
    end else begin
      if(io_deq_valid) begin
        if(GEN_49 == roq_deq_addr) begin
          roq_free_2 <= GEN_2;
        end else begin
          if(T_110) begin
            if(GEN_49 == roq_enq_addr) begin
              roq_free_2 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_110) begin
          if(GEN_49 == roq_enq_addr) begin
            roq_free_2 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_3 <= T_50_3;
    end else begin
      if(io_deq_valid) begin
        if(GEN_50 == roq_deq_addr) begin
          roq_free_3 <= GEN_2;
        end else begin
          if(T_110) begin
            if(GEN_50 == roq_enq_addr) begin
              roq_free_3 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_110) begin
          if(GEN_50 == roq_enq_addr) begin
            roq_free_3 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_4 <= T_50_4;
    end else begin
      if(io_deq_valid) begin
        if(3'h4 == roq_deq_addr) begin
          roq_free_4 <= GEN_2;
        end else begin
          if(T_110) begin
            if(3'h4 == roq_enq_addr) begin
              roq_free_4 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_110) begin
          if(3'h4 == roq_enq_addr) begin
            roq_free_4 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_5 <= T_50_5;
    end else begin
      if(io_deq_valid) begin
        if(3'h5 == roq_deq_addr) begin
          roq_free_5 <= GEN_2;
        end else begin
          if(T_110) begin
            if(3'h5 == roq_enq_addr) begin
              roq_free_5 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_110) begin
          if(3'h5 == roq_enq_addr) begin
            roq_free_5 <= GEN_1;
          end
        end
      end
    end
  end
endmodule
module ClientTileLinkIOUnwrapper(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [2:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_probe_ready,
  output  io_in_probe_valid,
  output [25:0] io_in_probe_bits_addr_block,
  output [1:0] io_in_probe_bits_p_type,
  output  io_in_release_ready,
  input   io_in_release_valid,
  input  [2:0] io_in_release_bits_addr_beat,
  input  [25:0] io_in_release_bits_addr_block,
  input  [2:0] io_in_release_bits_client_xact_id,
  input   io_in_release_bits_voluntary,
  input  [2:0] io_in_release_bits_r_type,
  input  [63:0] io_in_release_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [2:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  output  io_in_grant_bits_manager_id,
  output  io_in_finish_ready,
  input   io_in_finish_valid,
  input   io_in_finish_bits_manager_xact_id,
  input   io_in_finish_bits_manager_id,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  wire  acqArb_clk;
  wire  acqArb_reset;
  wire  acqArb_io_in_0_ready;
  wire  acqArb_io_in_0_valid;
  wire [25:0] acqArb_io_in_0_bits_addr_block;
  wire [2:0] acqArb_io_in_0_bits_client_xact_id;
  wire [2:0] acqArb_io_in_0_bits_addr_beat;
  wire  acqArb_io_in_0_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_0_bits_a_type;
  wire [11:0] acqArb_io_in_0_bits_union;
  wire [63:0] acqArb_io_in_0_bits_data;
  wire  acqArb_io_in_1_ready;
  wire  acqArb_io_in_1_valid;
  wire [25:0] acqArb_io_in_1_bits_addr_block;
  wire [2:0] acqArb_io_in_1_bits_client_xact_id;
  wire [2:0] acqArb_io_in_1_bits_addr_beat;
  wire  acqArb_io_in_1_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_1_bits_a_type;
  wire [11:0] acqArb_io_in_1_bits_union;
  wire [63:0] acqArb_io_in_1_bits_data;
  wire  acqArb_io_out_ready;
  wire  acqArb_io_out_valid;
  wire [25:0] acqArb_io_out_bits_addr_block;
  wire [2:0] acqArb_io_out_bits_client_xact_id;
  wire [2:0] acqArb_io_out_bits_addr_beat;
  wire  acqArb_io_out_bits_is_builtin_type;
  wire [2:0] acqArb_io_out_bits_a_type;
  wire [11:0] acqArb_io_out_bits_union;
  wire [63:0] acqArb_io_out_bits_data;
  wire  acqArb_io_chosen;
  wire  acqRoq_clk;
  wire  acqRoq_reset;
  wire  acqRoq_io_enq_ready;
  wire  acqRoq_io_enq_valid;
  wire  acqRoq_io_enq_bits_data;
  wire [2:0] acqRoq_io_enq_bits_tag;
  wire  acqRoq_io_deq_valid;
  wire [2:0] acqRoq_io_deq_tag;
  wire  acqRoq_io_deq_data;
  wire  acqRoq_io_deq_matches;
  wire  relRoq_clk;
  wire  relRoq_reset;
  wire  relRoq_io_enq_ready;
  wire  relRoq_io_enq_valid;
  wire  relRoq_io_enq_bits_data;
  wire [2:0] relRoq_io_enq_bits_tag;
  wire  relRoq_io_deq_valid;
  wire [2:0] relRoq_io_deq_tag;
  wire  relRoq_io_deq_data;
  wire  relRoq_io_deq_matches;
  wire [2:0] T_1366_0;
  wire  T_1368;
  wire  T_1371;
  wire  T_1373;
  wire [2:0] GEN_0;
  wire  T_1375;
  wire  acq_roq_enq;
  wire [2:0] T_1382_0;
  wire [2:0] T_1382_1;
  wire [2:0] T_1382_2;
  wire  T_1384;
  wire  T_1385;
  wire  T_1386;
  wire  T_1389;
  wire  T_1390;
  wire  T_1393;
  wire  T_1395;
  wire  rel_roq_enq;
  wire  T_1397;
  wire  acq_roq_ready;
  wire  T_1399;
  wire  rel_roq_ready;
  wire  T_1400;
  wire  T_1401;
  wire  T_1402;
  wire [2:0] T_1405;
  wire [11:0] T_1409;
  wire [25:0] T_1438_addr_block;
  wire [2:0] T_1438_client_xact_id;
  wire [2:0] T_1438_addr_beat;
  wire  T_1438_is_builtin_type;
  wire [2:0] T_1438_a_type;
  wire [11:0] T_1438_union;
  wire [63:0] T_1438_data;
  wire  T_1466;
  wire  T_1467;
  wire  T_1468;
  wire  T_1469;
  wire [7:0] GEN_2;
  wire [7:0] T_1493;
  wire [8:0] T_1538;
  wire [11:0] T_1556;
  wire [25:0] T_1591_addr_block;
  wire [2:0] T_1591_client_xact_id;
  wire [2:0] T_1591_addr_beat;
  wire  T_1591_is_builtin_type;
  wire [2:0] T_1591_a_type;
  wire [11:0] T_1591_union;
  wire [63:0] T_1591_data;
  wire  T_1619;
  wire  T_1620;
  wire [2:0] T_1628_0;
  wire [3:0] GEN_3;
  wire  T_1630;
  wire  T_1638_0;
  wire [3:0] GEN_4;
  wire  T_1640;
  wire  T_1643;
  wire  T_1646;
  wire  T_1648;
  wire  T_1649;
  wire  grant_deq_roq;
  wire  T_1650;
  wire  T_1652;
  wire  T_1653;
  wire  T_1655;
  wire  T_1656;
  wire  T_1657;
  wire  T_1658;
  wire  T_1660;
  wire [3:0] T_1661;
  wire [2:0] acq_grant_addr_beat;
  wire [2:0] acq_grant_client_xact_id;
  wire  acq_grant_manager_xact_id;
  wire  acq_grant_is_builtin_type;
  wire [3:0] acq_grant_g_type;
  wire [63:0] acq_grant_data;
  wire  T_1716;
  wire  T_1717;
  wire  T_1718;
  wire  T_1720;
  wire [2:0] rel_grant_addr_beat;
  wire [2:0] rel_grant_client_xact_id;
  wire  rel_grant_manager_xact_id;
  wire  rel_grant_is_builtin_type;
  wire [3:0] rel_grant_g_type;
  wire [63:0] rel_grant_data;
  wire [2:0] T_1776_addr_beat;
  wire [2:0] T_1776_client_xact_id;
  wire  T_1776_manager_xact_id;
  wire  T_1776_is_builtin_type;
  wire [3:0] T_1776_g_type;
  wire [63:0] T_1776_data;
  reg [25:0] GEN_1;
  reg [31:0] GEN_8;
  reg [1:0] GEN_5;
  reg [31:0] GEN_9;
  reg  GEN_6;
  reg [31:0] GEN_10;
  reg  GEN_7;
  reg [31:0] GEN_11;
  LockingRRArbiter_9 acqArb (
    .clk(acqArb_clk),
    .reset(acqArb_reset),
    .io_in_0_ready(acqArb_io_in_0_ready),
    .io_in_0_valid(acqArb_io_in_0_valid),
    .io_in_0_bits_addr_block(acqArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(acqArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(acqArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(acqArb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(acqArb_io_in_0_bits_a_type),
    .io_in_0_bits_union(acqArb_io_in_0_bits_union),
    .io_in_0_bits_data(acqArb_io_in_0_bits_data),
    .io_in_1_ready(acqArb_io_in_1_ready),
    .io_in_1_valid(acqArb_io_in_1_valid),
    .io_in_1_bits_addr_block(acqArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(acqArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(acqArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(acqArb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(acqArb_io_in_1_bits_a_type),
    .io_in_1_bits_union(acqArb_io_in_1_bits_union),
    .io_in_1_bits_data(acqArb_io_in_1_bits_data),
    .io_out_ready(acqArb_io_out_ready),
    .io_out_valid(acqArb_io_out_valid),
    .io_out_bits_addr_block(acqArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(acqArb_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(acqArb_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(acqArb_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(acqArb_io_out_bits_a_type),
    .io_out_bits_union(acqArb_io_out_bits_union),
    .io_out_bits_data(acqArb_io_out_bits_data),
    .io_chosen(acqArb_io_chosen)
  );
  ReorderQueue acqRoq (
    .clk(acqRoq_clk),
    .reset(acqRoq_reset),
    .io_enq_ready(acqRoq_io_enq_ready),
    .io_enq_valid(acqRoq_io_enq_valid),
    .io_enq_bits_data(acqRoq_io_enq_bits_data),
    .io_enq_bits_tag(acqRoq_io_enq_bits_tag),
    .io_deq_valid(acqRoq_io_deq_valid),
    .io_deq_tag(acqRoq_io_deq_tag),
    .io_deq_data(acqRoq_io_deq_data),
    .io_deq_matches(acqRoq_io_deq_matches)
  );
  ReorderQueue relRoq (
    .clk(relRoq_clk),
    .reset(relRoq_reset),
    .io_enq_ready(relRoq_io_enq_ready),
    .io_enq_valid(relRoq_io_enq_valid),
    .io_enq_bits_data(relRoq_io_enq_bits_data),
    .io_enq_bits_tag(relRoq_io_enq_bits_tag),
    .io_deq_valid(relRoq_io_deq_valid),
    .io_deq_tag(relRoq_io_deq_tag),
    .io_deq_data(relRoq_io_deq_data),
    .io_deq_matches(relRoq_io_deq_matches)
  );
  assign io_in_acquire_ready = T_1466;
  assign io_in_probe_valid = 1'h0;
  assign io_in_probe_bits_addr_block = GEN_1;
  assign io_in_probe_bits_p_type = GEN_5;
  assign io_in_release_ready = T_1619;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_grant_bits_addr_beat = T_1776_addr_beat;
  assign io_in_grant_bits_client_xact_id = T_1776_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = T_1776_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = T_1776_is_builtin_type;
  assign io_in_grant_bits_g_type = T_1776_g_type;
  assign io_in_grant_bits_data = T_1776_data;
  assign io_in_grant_bits_manager_id = GEN_6;
  assign io_in_finish_ready = GEN_7;
  assign io_out_acquire_valid = acqArb_io_out_valid;
  assign io_out_acquire_bits_addr_block = acqArb_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = acqArb_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = acqArb_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = acqArb_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = acqArb_io_out_bits_a_type;
  assign io_out_acquire_bits_union = acqArb_io_out_bits_union;
  assign io_out_acquire_bits_data = acqArb_io_out_bits_data;
  assign io_out_grant_ready = io_in_grant_ready;
  assign acqArb_clk = clk;
  assign acqArb_reset = reset;
  assign acqArb_io_in_0_valid = T_1402;
  assign acqArb_io_in_0_bits_addr_block = T_1438_addr_block;
  assign acqArb_io_in_0_bits_client_xact_id = T_1438_client_xact_id;
  assign acqArb_io_in_0_bits_addr_beat = T_1438_addr_beat;
  assign acqArb_io_in_0_bits_is_builtin_type = T_1438_is_builtin_type;
  assign acqArb_io_in_0_bits_a_type = T_1438_a_type;
  assign acqArb_io_in_0_bits_union = T_1438_union;
  assign acqArb_io_in_0_bits_data = T_1438_data;
  assign acqArb_io_in_1_valid = T_1469;
  assign acqArb_io_in_1_bits_addr_block = T_1591_addr_block;
  assign acqArb_io_in_1_bits_client_xact_id = T_1591_client_xact_id;
  assign acqArb_io_in_1_bits_addr_beat = T_1591_addr_beat;
  assign acqArb_io_in_1_bits_is_builtin_type = T_1591_is_builtin_type;
  assign acqArb_io_in_1_bits_a_type = T_1591_a_type;
  assign acqArb_io_in_1_bits_union = T_1591_union;
  assign acqArb_io_in_1_bits_data = T_1591_data;
  assign acqArb_io_out_ready = io_out_acquire_ready;
  assign acqRoq_clk = clk;
  assign acqRoq_reset = reset;
  assign acqRoq_io_enq_valid = T_1401;
  assign acqRoq_io_enq_bits_data = io_in_acquire_bits_is_builtin_type;
  assign acqRoq_io_enq_bits_tag = io_in_acquire_bits_client_xact_id;
  assign acqRoq_io_deq_valid = T_1650;
  assign acqRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign relRoq_clk = clk;
  assign relRoq_reset = reset;
  assign relRoq_io_enq_valid = T_1468;
  assign relRoq_io_enq_bits_data = io_in_release_bits_voluntary;
  assign relRoq_io_enq_bits_tag = io_in_release_bits_client_xact_id;
  assign relRoq_io_deq_valid = T_1653;
  assign relRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign T_1366_0 = 3'h3;
  assign T_1368 = T_1366_0 == io_in_acquire_bits_a_type;
  assign T_1371 = io_in_acquire_bits_is_builtin_type & T_1368;
  assign T_1373 = T_1371 == 1'h0;
  assign GEN_0 = {{2'd0}, 1'h0};
  assign T_1375 = io_in_acquire_bits_addr_beat == GEN_0;
  assign acq_roq_enq = T_1373 | T_1375;
  assign T_1382_0 = 3'h0;
  assign T_1382_1 = 3'h1;
  assign T_1382_2 = 3'h2;
  assign T_1384 = T_1382_0 == io_in_release_bits_r_type;
  assign T_1385 = T_1382_1 == io_in_release_bits_r_type;
  assign T_1386 = T_1382_2 == io_in_release_bits_r_type;
  assign T_1389 = T_1384 | T_1385;
  assign T_1390 = T_1389 | T_1386;
  assign T_1393 = T_1390 == 1'h0;
  assign T_1395 = io_in_release_bits_addr_beat == GEN_0;
  assign rel_roq_enq = T_1393 | T_1395;
  assign T_1397 = acq_roq_enq == 1'h0;
  assign acq_roq_ready = T_1397 | acqRoq_io_enq_ready;
  assign T_1399 = rel_roq_enq == 1'h0;
  assign rel_roq_ready = T_1399 | relRoq_io_enq_ready;
  assign T_1400 = io_in_acquire_valid & acqArb_io_in_0_ready;
  assign T_1401 = T_1400 & acq_roq_enq;
  assign T_1402 = io_in_acquire_valid & acq_roq_ready;
  assign T_1405 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_a_type : 3'h1;
  assign T_1409 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_union : {{3'd0}, 9'h1c1};
  assign T_1438_addr_block = io_in_acquire_bits_addr_block;
  assign T_1438_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign T_1438_addr_beat = io_in_acquire_bits_addr_beat;
  assign T_1438_is_builtin_type = 1'h1;
  assign T_1438_a_type = T_1405;
  assign T_1438_union = T_1409;
  assign T_1438_data = io_in_acquire_bits_data;
  assign T_1466 = acq_roq_ready & acqArb_io_in_0_ready;
  assign T_1467 = io_in_release_valid & acqArb_io_in_1_ready;
  assign T_1468 = T_1467 & rel_roq_enq;
  assign T_1469 = io_in_release_valid & rel_roq_ready;
  assign GEN_2 = $signed(8'hff);
  assign T_1493 = $unsigned(GEN_2);
  assign T_1538 = {T_1493,1'h1};
  assign T_1556 = 1'h1 ? {{3'd0}, T_1538} : 12'h0;
  assign T_1591_addr_block = io_in_release_bits_addr_block;
  assign T_1591_client_xact_id = io_in_release_bits_client_xact_id;
  assign T_1591_addr_beat = io_in_release_bits_addr_beat;
  assign T_1591_is_builtin_type = 1'h1;
  assign T_1591_a_type = 3'h3;
  assign T_1591_union = T_1556;
  assign T_1591_data = io_in_release_bits_data;
  assign T_1619 = rel_roq_ready & acqArb_io_in_1_ready;
  assign T_1620 = io_out_grant_ready & io_out_grant_valid;
  assign T_1628_0 = 3'h5;
  assign GEN_3 = {{1'd0}, T_1628_0};
  assign T_1630 = GEN_3 == io_out_grant_bits_g_type;
  assign T_1638_0 = 1'h0;
  assign GEN_4 = {{3'd0}, T_1638_0};
  assign T_1640 = GEN_4 == io_out_grant_bits_g_type;
  assign T_1643 = io_out_grant_bits_is_builtin_type ? T_1630 : T_1640;
  assign T_1646 = T_1643 == 1'h0;
  assign T_1648 = io_out_grant_bits_addr_beat == 3'h7;
  assign T_1649 = T_1646 | T_1648;
  assign grant_deq_roq = T_1620 & T_1649;
  assign T_1650 = acqRoq_io_deq_matches & grant_deq_roq;
  assign T_1652 = acqRoq_io_deq_matches == 1'h0;
  assign T_1653 = T_1652 & grant_deq_roq;
  assign T_1655 = grant_deq_roq == 1'h0;
  assign T_1656 = T_1655 | acqRoq_io_deq_matches;
  assign T_1657 = T_1656 | relRoq_io_deq_matches;
  assign T_1658 = T_1657 | reset;
  assign T_1660 = T_1658 == 1'h0;
  assign T_1661 = acqRoq_io_deq_data ? io_out_grant_bits_g_type : {{3'd0}, 1'h0};
  assign acq_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign acq_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign acq_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign acq_grant_is_builtin_type = acqRoq_io_deq_data;
  assign acq_grant_g_type = T_1661;
  assign acq_grant_data = io_out_grant_bits_data;
  assign T_1716 = io_in_release_valid == 1'h0;
  assign T_1717 = T_1716 | io_in_release_bits_voluntary;
  assign T_1718 = T_1717 | reset;
  assign T_1720 = T_1718 == 1'h0;
  assign rel_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign rel_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign rel_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign rel_grant_is_builtin_type = 1'h1;
  assign rel_grant_g_type = {{1'd0}, 3'h0};
  assign rel_grant_data = io_out_grant_bits_data;
  assign T_1776_addr_beat = acqRoq_io_deq_matches ? acq_grant_addr_beat : rel_grant_addr_beat;
  assign T_1776_client_xact_id = acqRoq_io_deq_matches ? acq_grant_client_xact_id : rel_grant_client_xact_id;
  assign T_1776_manager_xact_id = acqRoq_io_deq_matches ? acq_grant_manager_xact_id : rel_grant_manager_xact_id;
  assign T_1776_is_builtin_type = acqRoq_io_deq_matches ? acq_grant_is_builtin_type : rel_grant_is_builtin_type;
  assign T_1776_g_type = acqRoq_io_deq_matches ? acq_grant_g_type : rel_grant_g_type;
  assign T_1776_data = acqRoq_io_deq_matches ? acq_grant_data : rel_grant_data;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_8 = {1{$random}};
  GEN_1 = GEN_8[25:0];
  GEN_9 = {1{$random}};
  GEN_5 = GEN_9[1:0];
  GEN_10 = {1{$random}};
  GEN_6 = GEN_10[0:0];
  GEN_11 = {1{$random}};
  GEN_7 = GEN_11[0:0];
  end
`endif
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1660) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink Unwrapper: client_xact_id mismatch\n    at Tilelink.scala:123 assert(!grant_deq_roq || acqRoq.io.deq.matches || relRoq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1660) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1660) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1720) begin
          $fwrite(32'h80000002,"Assertion failed: Unwrapper can only process voluntary releases.\n    at Tilelink.scala:137 assert(!io.in.release.valid || io.in.release.bits.isVoluntary(), \"Unwrapper can only process voluntary releases.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1720) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1720) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientTileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [2:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [2:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [2:0] io_inner_grant_bits_client_xact_id,
  output  io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_manager_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input   io_inner_finish_bits_manager_xact_id,
  input   io_inner_finish_bits_manager_id,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  assign io_inner_acquire_ready = io_outer_acquire_ready;
  assign io_inner_probe_valid = io_outer_probe_valid;
  assign io_inner_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign io_inner_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign io_inner_release_ready = io_outer_release_ready;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_manager_id = io_outer_grant_bits_manager_id;
  assign io_inner_finish_ready = io_outer_finish_ready;
  assign io_outer_acquire_valid = io_inner_acquire_valid;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_probe_ready = io_inner_probe_ready;
  assign io_outer_release_valid = io_inner_release_valid;
  assign io_outer_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign io_outer_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign io_outer_release_bits_r_type = io_inner_release_bits_r_type;
  assign io_outer_release_bits_data = io_inner_release_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_finish_valid = io_inner_finish_valid;
  assign io_outer_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign io_outer_finish_bits_manager_id = io_inner_finish_bits_manager_id;
endmodule
module ReorderQueue_2(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_data_addr_beat,
  input   io_enq_bits_data_subblock,
  input  [4:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [4:0] io_deq_tag,
  output [2:0] io_deq_data_addr_beat,
  output  io_deq_data_subblock,
  output  io_deq_matches
);
  reg [2:0] roq_data_addr_beat [0:5];
  reg [31:0] GEN_15;
  wire [2:0] roq_data_addr_beat_T_324_data;
  wire [2:0] roq_data_addr_beat_T_324_addr;
  wire  roq_data_addr_beat_T_324_en;
  wire [2:0] roq_data_addr_beat_T_353_data;
  wire [2:0] roq_data_addr_beat_T_353_addr;
  wire  roq_data_addr_beat_T_353_mask;
  wire  roq_data_addr_beat_T_353_en;
  reg  roq_data_subblock [0:5];
  reg [31:0] GEN_16;
  wire  roq_data_subblock_T_324_data;
  wire [2:0] roq_data_subblock_T_324_addr;
  wire  roq_data_subblock_T_324_en;
  wire  roq_data_subblock_T_353_data;
  wire [2:0] roq_data_subblock_T_353_addr;
  wire  roq_data_subblock_T_353_mask;
  wire  roq_data_subblock_T_353_en;
  reg [4:0] roq_tags_0;
  reg [31:0] GEN_17;
  reg [4:0] roq_tags_1;
  reg [31:0] GEN_18;
  reg [4:0] roq_tags_2;
  reg [31:0] GEN_19;
  reg [4:0] roq_tags_3;
  reg [31:0] GEN_20;
  reg [4:0] roq_tags_4;
  reg [31:0] GEN_21;
  reg [4:0] roq_tags_5;
  reg [31:0] GEN_22;
  wire  T_270_0;
  wire  T_270_1;
  wire  T_270_2;
  wire  T_270_3;
  wire  T_270_4;
  wire  T_270_5;
  reg  roq_free_0;
  reg [31:0] GEN_29;
  reg  roq_free_1;
  reg [31:0] GEN_42;
  reg  roq_free_2;
  reg [31:0] GEN_53;
  reg  roq_free_3;
  reg [31:0] GEN_54;
  reg  roq_free_4;
  reg [31:0] GEN_55;
  reg  roq_free_5;
  reg [31:0] GEN_56;
  wire [2:0] T_281;
  wire [2:0] T_282;
  wire [2:0] T_283;
  wire [2:0] T_284;
  wire [2:0] roq_enq_addr;
  wire  T_285;
  wire  T_287;
  wire  T_288;
  wire  T_289;
  wire  T_291;
  wire  T_292;
  wire  T_293;
  wire  T_295;
  wire  T_296;
  wire  T_297;
  wire  T_299;
  wire  T_300;
  wire  T_301;
  wire  T_303;
  wire  T_304;
  wire  T_305;
  wire  T_307;
  wire  T_308;
  wire [2:0] T_315;
  wire [2:0] T_316;
  wire [2:0] T_317;
  wire [2:0] T_318;
  wire [2:0] roq_deq_addr;
  wire  T_319;
  wire  T_320;
  wire  T_321;
  wire  T_322;
  wire  T_323;
  wire  T_347;
  wire  T_348;
  wire  T_349;
  wire  T_350;
  wire  T_351;
  wire  T_352;
  wire [4:0] GEN_0;
  wire [2:0] GEN_49;
  wire [4:0] GEN_3;
  wire [2:0] GEN_50;
  wire [4:0] GEN_4;
  wire [2:0] GEN_51;
  wire [4:0] GEN_5;
  wire [2:0] GEN_52;
  wire [4:0] GEN_6;
  wire [4:0] GEN_7;
  wire [4:0] GEN_8;
  wire  GEN_1;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [4:0] GEN_23;
  wire [4:0] GEN_24;
  wire [4:0] GEN_25;
  wire [4:0] GEN_26;
  wire [4:0] GEN_27;
  wire [4:0] GEN_28;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_2;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  assign io_enq_ready = T_323;
  assign io_deq_data_addr_beat = roq_data_addr_beat_T_324_data;
  assign io_deq_data_subblock = roq_data_subblock_T_324_data;
  assign io_deq_matches = T_351;
  assign roq_data_addr_beat_T_324_addr = roq_deq_addr;
  assign roq_data_addr_beat_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_addr_beat_T_324_data = roq_data_addr_beat[roq_data_addr_beat_T_324_addr];
  `else
  assign roq_data_addr_beat_T_324_data = roq_data_addr_beat_T_324_addr >= 3'h6 ? $random : roq_data_addr_beat[roq_data_addr_beat_T_324_addr];
  `endif
  assign roq_data_addr_beat_T_353_data = io_enq_bits_data_addr_beat;
  assign roq_data_addr_beat_T_353_addr = roq_enq_addr;
  assign roq_data_addr_beat_T_353_mask = T_352;
  assign roq_data_addr_beat_T_353_en = T_352;
  assign roq_data_subblock_T_324_addr = roq_deq_addr;
  assign roq_data_subblock_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_subblock_T_324_data = roq_data_subblock[roq_data_subblock_T_324_addr];
  `else
  assign roq_data_subblock_T_324_data = roq_data_subblock_T_324_addr >= 3'h6 ? $random : roq_data_subblock[roq_data_subblock_T_324_addr];
  `endif
  assign roq_data_subblock_T_353_data = io_enq_bits_data_subblock;
  assign roq_data_subblock_T_353_addr = roq_enq_addr;
  assign roq_data_subblock_T_353_mask = T_352;
  assign roq_data_subblock_T_353_en = T_352;
  assign T_270_0 = 1'h1;
  assign T_270_1 = 1'h1;
  assign T_270_2 = 1'h1;
  assign T_270_3 = 1'h1;
  assign T_270_4 = 1'h1;
  assign T_270_5 = 1'h1;
  assign T_281 = roq_free_4 ? 3'h4 : 3'h5;
  assign T_282 = roq_free_3 ? {{1'd0}, 2'h3} : T_281;
  assign T_283 = roq_free_2 ? {{1'd0}, 2'h2} : T_282;
  assign T_284 = roq_free_1 ? {{2'd0}, 1'h1} : T_283;
  assign roq_enq_addr = roq_free_0 ? {{2'd0}, 1'h0} : T_284;
  assign T_285 = roq_tags_0 == io_deq_tag;
  assign T_287 = roq_free_0 == 1'h0;
  assign T_288 = T_285 & T_287;
  assign T_289 = roq_tags_1 == io_deq_tag;
  assign T_291 = roq_free_1 == 1'h0;
  assign T_292 = T_289 & T_291;
  assign T_293 = roq_tags_2 == io_deq_tag;
  assign T_295 = roq_free_2 == 1'h0;
  assign T_296 = T_293 & T_295;
  assign T_297 = roq_tags_3 == io_deq_tag;
  assign T_299 = roq_free_3 == 1'h0;
  assign T_300 = T_297 & T_299;
  assign T_301 = roq_tags_4 == io_deq_tag;
  assign T_303 = roq_free_4 == 1'h0;
  assign T_304 = T_301 & T_303;
  assign T_305 = roq_tags_5 == io_deq_tag;
  assign T_307 = roq_free_5 == 1'h0;
  assign T_308 = T_305 & T_307;
  assign T_315 = T_304 ? 3'h4 : 3'h5;
  assign T_316 = T_300 ? {{1'd0}, 2'h3} : T_315;
  assign T_317 = T_296 ? {{1'd0}, 2'h2} : T_316;
  assign T_318 = T_292 ? {{2'd0}, 1'h1} : T_317;
  assign roq_deq_addr = T_288 ? {{2'd0}, 1'h0} : T_318;
  assign T_319 = roq_free_0 | roq_free_1;
  assign T_320 = T_319 | roq_free_2;
  assign T_321 = T_320 | roq_free_3;
  assign T_322 = T_321 | roq_free_4;
  assign T_323 = T_322 | roq_free_5;
  assign T_347 = T_288 | T_292;
  assign T_348 = T_347 | T_296;
  assign T_349 = T_348 | T_300;
  assign T_350 = T_349 | T_304;
  assign T_351 = T_350 | T_308;
  assign T_352 = io_enq_valid & io_enq_ready;
  assign GEN_0 = io_enq_bits_tag;
  assign GEN_49 = {{2'd0}, 1'h0};
  assign GEN_3 = GEN_49 == roq_enq_addr ? GEN_0 : roq_tags_0;
  assign GEN_50 = {{2'd0}, 1'h1};
  assign GEN_4 = GEN_50 == roq_enq_addr ? GEN_0 : roq_tags_1;
  assign GEN_51 = {{1'd0}, 2'h2};
  assign GEN_5 = GEN_51 == roq_enq_addr ? GEN_0 : roq_tags_2;
  assign GEN_52 = {{1'd0}, 2'h3};
  assign GEN_6 = GEN_52 == roq_enq_addr ? GEN_0 : roq_tags_3;
  assign GEN_7 = 3'h4 == roq_enq_addr ? GEN_0 : roq_tags_4;
  assign GEN_8 = 3'h5 == roq_enq_addr ? GEN_0 : roq_tags_5;
  assign GEN_1 = 1'h0;
  assign GEN_9 = GEN_49 == roq_enq_addr ? GEN_1 : roq_free_0;
  assign GEN_10 = GEN_50 == roq_enq_addr ? GEN_1 : roq_free_1;
  assign GEN_11 = GEN_51 == roq_enq_addr ? GEN_1 : roq_free_2;
  assign GEN_12 = GEN_52 == roq_enq_addr ? GEN_1 : roq_free_3;
  assign GEN_13 = 3'h4 == roq_enq_addr ? GEN_1 : roq_free_4;
  assign GEN_14 = 3'h5 == roq_enq_addr ? GEN_1 : roq_free_5;
  assign GEN_23 = T_352 ? GEN_3 : roq_tags_0;
  assign GEN_24 = T_352 ? GEN_4 : roq_tags_1;
  assign GEN_25 = T_352 ? GEN_5 : roq_tags_2;
  assign GEN_26 = T_352 ? GEN_6 : roq_tags_3;
  assign GEN_27 = T_352 ? GEN_7 : roq_tags_4;
  assign GEN_28 = T_352 ? GEN_8 : roq_tags_5;
  assign GEN_30 = T_352 ? GEN_9 : roq_free_0;
  assign GEN_31 = T_352 ? GEN_10 : roq_free_1;
  assign GEN_32 = T_352 ? GEN_11 : roq_free_2;
  assign GEN_33 = T_352 ? GEN_12 : roq_free_3;
  assign GEN_34 = T_352 ? GEN_13 : roq_free_4;
  assign GEN_35 = T_352 ? GEN_14 : roq_free_5;
  assign GEN_2 = 1'h1;
  assign GEN_36 = GEN_49 == roq_deq_addr ? GEN_2 : GEN_30;
  assign GEN_37 = GEN_50 == roq_deq_addr ? GEN_2 : GEN_31;
  assign GEN_38 = GEN_51 == roq_deq_addr ? GEN_2 : GEN_32;
  assign GEN_39 = GEN_52 == roq_deq_addr ? GEN_2 : GEN_33;
  assign GEN_40 = 3'h4 == roq_deq_addr ? GEN_2 : GEN_34;
  assign GEN_41 = 3'h5 == roq_deq_addr ? GEN_2 : GEN_35;
  assign GEN_43 = io_deq_valid ? GEN_36 : GEN_30;
  assign GEN_44 = io_deq_valid ? GEN_37 : GEN_31;
  assign GEN_45 = io_deq_valid ? GEN_38 : GEN_32;
  assign GEN_46 = io_deq_valid ? GEN_39 : GEN_33;
  assign GEN_47 = io_deq_valid ? GEN_40 : GEN_34;
  assign GEN_48 = io_deq_valid ? GEN_41 : GEN_35;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    roq_data_addr_beat[initvar] = GEN_15[2:0];
  GEN_16 = {1{$random}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    roq_data_subblock[initvar] = GEN_16[0:0];
  GEN_17 = {1{$random}};
  roq_tags_0 = GEN_17[4:0];
  GEN_18 = {1{$random}};
  roq_tags_1 = GEN_18[4:0];
  GEN_19 = {1{$random}};
  roq_tags_2 = GEN_19[4:0];
  GEN_20 = {1{$random}};
  roq_tags_3 = GEN_20[4:0];
  GEN_21 = {1{$random}};
  roq_tags_4 = GEN_21[4:0];
  GEN_22 = {1{$random}};
  roq_tags_5 = GEN_22[4:0];
  GEN_29 = {1{$random}};
  roq_free_0 = GEN_29[0:0];
  GEN_42 = {1{$random}};
  roq_free_1 = GEN_42[0:0];
  GEN_53 = {1{$random}};
  roq_free_2 = GEN_53[0:0];
  GEN_54 = {1{$random}};
  roq_free_3 = GEN_54[0:0];
  GEN_55 = {1{$random}};
  roq_free_4 = GEN_55[0:0];
  GEN_56 = {1{$random}};
  roq_free_5 = GEN_56[0:0];
  end
`endif
  always @(posedge clk) begin
    if(roq_data_addr_beat_T_353_en & roq_data_addr_beat_T_353_mask) begin
      roq_data_addr_beat[roq_data_addr_beat_T_353_addr] <= roq_data_addr_beat_T_353_data;
    end
    if(roq_data_subblock_T_353_en & roq_data_subblock_T_353_mask) begin
      roq_data_subblock[roq_data_subblock_T_353_addr] <= roq_data_subblock_T_353_data;
    end
    if(1'h0) begin
    end else begin
      if(T_352) begin
        if(GEN_49 == roq_enq_addr) begin
          roq_tags_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_352) begin
        if(GEN_50 == roq_enq_addr) begin
          roq_tags_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_352) begin
        if(GEN_51 == roq_enq_addr) begin
          roq_tags_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_352) begin
        if(GEN_52 == roq_enq_addr) begin
          roq_tags_3 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_352) begin
        if(3'h4 == roq_enq_addr) begin
          roq_tags_4 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_352) begin
        if(3'h5 == roq_enq_addr) begin
          roq_tags_5 <= GEN_0;
        end
      end
    end
    if(reset) begin
      roq_free_0 <= T_270_0;
    end else begin
      if(io_deq_valid) begin
        if(GEN_49 == roq_deq_addr) begin
          roq_free_0 <= GEN_2;
        end else begin
          if(T_352) begin
            if(GEN_49 == roq_enq_addr) begin
              roq_free_0 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_352) begin
          if(GEN_49 == roq_enq_addr) begin
            roq_free_0 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_1 <= T_270_1;
    end else begin
      if(io_deq_valid) begin
        if(GEN_50 == roq_deq_addr) begin
          roq_free_1 <= GEN_2;
        end else begin
          if(T_352) begin
            if(GEN_50 == roq_enq_addr) begin
              roq_free_1 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_352) begin
          if(GEN_50 == roq_enq_addr) begin
            roq_free_1 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_2 <= T_270_2;
    end else begin
      if(io_deq_valid) begin
        if(GEN_51 == roq_deq_addr) begin
          roq_free_2 <= GEN_2;
        end else begin
          if(T_352) begin
            if(GEN_51 == roq_enq_addr) begin
              roq_free_2 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_352) begin
          if(GEN_51 == roq_enq_addr) begin
            roq_free_2 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_3 <= T_270_3;
    end else begin
      if(io_deq_valid) begin
        if(GEN_52 == roq_deq_addr) begin
          roq_free_3 <= GEN_2;
        end else begin
          if(T_352) begin
            if(GEN_52 == roq_enq_addr) begin
              roq_free_3 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_352) begin
          if(GEN_52 == roq_enq_addr) begin
            roq_free_3 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_4 <= T_270_4;
    end else begin
      if(io_deq_valid) begin
        if(3'h4 == roq_deq_addr) begin
          roq_free_4 <= GEN_2;
        end else begin
          if(T_352) begin
            if(3'h4 == roq_enq_addr) begin
              roq_free_4 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_352) begin
          if(3'h4 == roq_enq_addr) begin
            roq_free_4 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_5 <= T_270_5;
    end else begin
      if(io_deq_valid) begin
        if(3'h5 == roq_deq_addr) begin
          roq_free_5 <= GEN_2;
        end else begin
          if(T_352) begin
            if(3'h5 == roq_enq_addr) begin
              roq_free_5 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_352) begin
          if(3'h5 == roq_enq_addr) begin
            roq_free_5 <= GEN_1;
          end
        end
      end
    end
  end
endmodule
module NastiIOTileLinkIOIdMapper(
  input   clk,
  input   reset,
  input   io_req_valid,
  output  io_req_ready,
  input  [2:0] io_req_tl_id,
  output [4:0] io_req_nasti_id,
  input   io_resp_valid,
  output  io_resp_matches,
  input  [4:0] io_resp_nasti_id,
  output [2:0] io_resp_tl_id
);
  assign io_req_ready = 1'h1;
  assign io_req_nasti_id = {{2'd0}, io_req_tl_id};
  assign io_resp_matches = 1'h1;
  assign io_resp_tl_id = io_resp_nasti_id[2:0];
endmodule
module Arbiter_13(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [2:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [2:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [2:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output  io_chosen
);
  wire  GEN_0;
  wire [2:0] GEN_1;
  wire [2:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire [3:0] GEN_5;
  wire [63:0] GEN_6;
  wire  GEN_7;
  wire  T_652;
  wire  T_654;
  wire  T_656;
  wire  T_657;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_654;
  assign io_out_valid = T_657;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_client_id = GEN_7;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr_beat : io_in_1_bits_addr_beat;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_client_xact_id : io_in_1_bits_client_xact_id;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_manager_xact_id : io_in_1_bits_manager_xact_id;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_is_builtin_type : io_in_1_bits_is_builtin_type;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_g_type : io_in_1_bits_g_type;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_client_id : io_in_1_bits_client_id;
  assign T_652 = io_in_0_valid == 1'h0;
  assign T_654 = T_652 & io_out_ready;
  assign T_656 = T_652 == 1'h0;
  assign T_657 = T_656 | io_in_1_valid;
endmodule
module NastiIOTileLinkIOConverter(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [2:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [2:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  input   io_nasti_aw_ready,
  output  io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  output [7:0] io_nasti_aw_bits_len,
  output [2:0] io_nasti_aw_bits_size,
  output [1:0] io_nasti_aw_bits_burst,
  output  io_nasti_aw_bits_lock,
  output [3:0] io_nasti_aw_bits_cache,
  output [2:0] io_nasti_aw_bits_prot,
  output [3:0] io_nasti_aw_bits_qos,
  output [3:0] io_nasti_aw_bits_region,
  output [4:0] io_nasti_aw_bits_id,
  output  io_nasti_aw_bits_user,
  input   io_nasti_w_ready,
  output  io_nasti_w_valid,
  output [63:0] io_nasti_w_bits_data,
  output  io_nasti_w_bits_last,
  output [4:0] io_nasti_w_bits_id,
  output [7:0] io_nasti_w_bits_strb,
  output  io_nasti_w_bits_user,
  output  io_nasti_b_ready,
  input   io_nasti_b_valid,
  input  [1:0] io_nasti_b_bits_resp,
  input  [4:0] io_nasti_b_bits_id,
  input   io_nasti_b_bits_user,
  input   io_nasti_ar_ready,
  output  io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output [7:0] io_nasti_ar_bits_len,
  output [2:0] io_nasti_ar_bits_size,
  output [1:0] io_nasti_ar_bits_burst,
  output  io_nasti_ar_bits_lock,
  output [3:0] io_nasti_ar_bits_cache,
  output [2:0] io_nasti_ar_bits_prot,
  output [3:0] io_nasti_ar_bits_qos,
  output [3:0] io_nasti_ar_bits_region,
  output [4:0] io_nasti_ar_bits_id,
  output  io_nasti_ar_bits_user,
  output  io_nasti_r_ready,
  input   io_nasti_r_valid,
  input  [1:0] io_nasti_r_bits_resp,
  input  [63:0] io_nasti_r_bits_data,
  input   io_nasti_r_bits_last,
  input  [4:0] io_nasti_r_bits_id,
  input   io_nasti_r_bits_user
);
  wire [2:0] T_688_0;
  wire [2:0] T_688_1;
  wire [2:0] T_688_2;
  wire  T_690;
  wire  T_691;
  wire  T_692;
  wire  T_695;
  wire  T_696;
  wire  has_data;
  wire [2:0] T_705_0;
  wire [2:0] T_705_1;
  wire [2:0] T_705_2;
  wire  T_707;
  wire  T_708;
  wire  T_709;
  wire  T_712;
  wire  T_713;
  wire  is_subblock;
  wire [2:0] T_722_0;
  wire  T_724;
  wire  is_multibeat;
  wire  T_727;
  wire  T_728;
  reg [2:0] tl_cnt_out;
  reg [31:0] GEN_15;
  wire  T_731;
  wire [2:0] GEN_6;
  wire [3:0] T_733;
  wire [2:0] T_734;
  wire [2:0] GEN_0;
  wire  tl_wrap_out;
  wire  T_736;
  wire  get_valid;
  wire  put_valid;
  wire  roq_clk;
  wire  roq_reset;
  wire  roq_io_enq_ready;
  wire  roq_io_enq_valid;
  wire [2:0] roq_io_enq_bits_data_addr_beat;
  wire  roq_io_enq_bits_data_subblock;
  wire [4:0] roq_io_enq_bits_tag;
  wire  roq_io_deq_valid;
  wire [4:0] roq_io_deq_tag;
  wire [2:0] roq_io_deq_data_addr_beat;
  wire  roq_io_deq_data_subblock;
  wire  roq_io_deq_matches;
  wire  get_id_mapper_clk;
  wire  get_id_mapper_reset;
  wire  get_id_mapper_io_req_valid;
  wire  get_id_mapper_io_req_ready;
  wire [2:0] get_id_mapper_io_req_tl_id;
  wire [4:0] get_id_mapper_io_req_nasti_id;
  wire  get_id_mapper_io_resp_valid;
  wire  get_id_mapper_io_resp_matches;
  wire [4:0] get_id_mapper_io_resp_nasti_id;
  wire [2:0] get_id_mapper_io_resp_tl_id;
  wire  put_id_mapper_clk;
  wire  put_id_mapper_reset;
  wire  put_id_mapper_io_req_valid;
  wire  put_id_mapper_io_req_ready;
  wire [2:0] put_id_mapper_io_req_tl_id;
  wire [4:0] put_id_mapper_io_req_nasti_id;
  wire  put_id_mapper_io_resp_valid;
  wire  put_id_mapper_io_resp_matches;
  wire [4:0] put_id_mapper_io_resp_nasti_id;
  wire [2:0] put_id_mapper_io_resp_tl_id;
  wire [2:0] GEN_7;
  wire  T_761;
  wire  put_id_mask;
  wire  T_763;
  wire  put_id_ready;
  reg  w_inflight;
  reg [31:0] GEN_16;
  wire  aw_ready;
  wire  T_765;
  wire  T_767;
  wire  T_768;
  reg [2:0] nasti_cnt_out;
  reg [31:0] GEN_17;
  wire  T_771;
  wire [3:0] T_773;
  wire [2:0] T_774;
  wire [2:0] GEN_1;
  wire  nasti_wrap_out;
  wire  T_775;
  wire  T_776;
  wire  T_778;
  wire  T_779;
  wire  T_780;
  wire  T_781;
  wire  T_783;
  wire  T_784;
  wire  T_785;
  wire  T_786;
  wire  T_787;
  wire  T_789;
  wire [2:0] T_790;
  wire [28:0] T_791;
  wire [31:0] T_792;
  wire [2:0] T_793;
  wire  T_803;
  wire [2:0] T_804;
  wire  T_805;
  wire [2:0] T_806;
  wire  T_807;
  wire [2:0] T_808;
  wire  T_809;
  wire [2:0] T_810;
  wire  T_811;
  wire [2:0] T_812;
  wire  T_813;
  wire [2:0] T_814;
  wire  T_815;
  wire [2:0] T_816;
  wire  T_817;
  wire [2:0] T_818;
  wire [2:0] T_820;
  wire [2:0] T_823;
  wire [31:0] T_843_addr;
  wire [7:0] T_843_len;
  wire [2:0] T_843_size;
  wire [1:0] T_843_burst;
  wire  T_843_lock;
  wire [3:0] T_843_cache;
  wire [2:0] T_843_prot;
  wire [3:0] T_843_qos;
  wire [3:0] T_843_region;
  wire [4:0] T_843_id;
  wire  T_843_user;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire  T_865;
  wire [2:0] T_872;
  wire [31:0] T_885_addr;
  wire [7:0] T_885_len;
  wire [2:0] T_885_size;
  wire [1:0] T_885_burst;
  wire  T_885_lock;
  wire [3:0] T_885_cache;
  wire [2:0] T_885_prot;
  wire [3:0] T_885_qos;
  wire [3:0] T_885_region;
  wire [4:0] T_885_id;
  wire  T_885_user;
  wire  T_904;
  wire  T_906;
  wire  T_907;
  wire [7:0] GEN_9;
  wire [8:0] T_911;
  wire [7:0] T_912;
  wire [7:0] T_918_0;
  wire  T_921;
  wire  T_922;
  wire  T_924;
  wire  T_925;
  wire  T_926;
  wire [7:0] T_927;
  wire [7:0] T_929;
  wire [7:0] T_930;
  wire  T_932;
  wire  T_933;
  wire [63:0] T_940_data;
  wire  T_940_last;
  wire [4:0] T_940_id;
  wire [7:0] T_940_strb;
  wire  T_940_user;
  wire  T_951;
  wire  T_952;
  wire  T_953;
  wire  T_954;
  wire  T_955;
  wire  T_959;
  wire  T_960;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  T_963;
  wire [2:0] T_971_0;
  wire [3:0] GEN_10;
  wire  T_973;
  wire  T_981_0;
  wire [3:0] GEN_11;
  wire  T_983;
  wire  T_986;
  wire  T_988;
  reg [2:0] tl_cnt_in;
  reg [31:0] GEN_18;
  wire [3:0] T_993;
  wire [2:0] T_994;
  wire [2:0] GEN_5;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [2:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_0_bits_client_id;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [2:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_1_bits_client_id;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [2:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_out_bits_client_id;
  wire  gnt_arb_io_chosen;
  wire [2:0] T_1026;
  wire [2:0] T_1028;
  wire [2:0] T_1056_addr_beat;
  wire [2:0] T_1056_client_xact_id;
  wire  T_1056_manager_xact_id;
  wire  T_1056_is_builtin_type;
  wire [3:0] T_1056_g_type;
  wire [63:0] T_1056_data;
  wire  T_1084;
  wire  T_1085;
  wire  T_1086;
  wire  T_1088;
  wire  T_1090;
  wire  T_1091;
  wire  T_1092;
  wire  T_1094;
  wire [2:0] T_1127_addr_beat;
  wire [2:0] T_1127_client_xact_id;
  wire  T_1127_manager_xact_id;
  wire  T_1127_is_builtin_type;
  wire [3:0] T_1127_g_type;
  wire [63:0] T_1127_data;
  wire  T_1155;
  wire  T_1156;
  wire  T_1157;
  wire  T_1159;
  wire  T_1161;
  wire [1:0] GEN_13;
  wire  T_1163;
  wire  T_1164;
  wire  T_1165;
  wire  T_1167;
  wire  T_1169;
  wire  T_1171;
  wire  T_1172;
  wire  T_1173;
  wire  T_1175;
  reg [4:0] GEN_8;
  reg [31:0] GEN_19;
  reg  GEN_12;
  reg [31:0] GEN_20;
  reg  GEN_14;
  reg [31:0] GEN_21;
  ReorderQueue_2 roq (
    .clk(roq_clk),
    .reset(roq_reset),
    .io_enq_ready(roq_io_enq_ready),
    .io_enq_valid(roq_io_enq_valid),
    .io_enq_bits_data_addr_beat(roq_io_enq_bits_data_addr_beat),
    .io_enq_bits_data_subblock(roq_io_enq_bits_data_subblock),
    .io_enq_bits_tag(roq_io_enq_bits_tag),
    .io_deq_valid(roq_io_deq_valid),
    .io_deq_tag(roq_io_deq_tag),
    .io_deq_data_addr_beat(roq_io_deq_data_addr_beat),
    .io_deq_data_subblock(roq_io_deq_data_subblock),
    .io_deq_matches(roq_io_deq_matches)
  );
  NastiIOTileLinkIOIdMapper get_id_mapper (
    .clk(get_id_mapper_clk),
    .reset(get_id_mapper_reset),
    .io_req_valid(get_id_mapper_io_req_valid),
    .io_req_ready(get_id_mapper_io_req_ready),
    .io_req_tl_id(get_id_mapper_io_req_tl_id),
    .io_req_nasti_id(get_id_mapper_io_req_nasti_id),
    .io_resp_valid(get_id_mapper_io_resp_valid),
    .io_resp_matches(get_id_mapper_io_resp_matches),
    .io_resp_nasti_id(get_id_mapper_io_resp_nasti_id),
    .io_resp_tl_id(get_id_mapper_io_resp_tl_id)
  );
  NastiIOTileLinkIOIdMapper put_id_mapper (
    .clk(put_id_mapper_clk),
    .reset(put_id_mapper_reset),
    .io_req_valid(put_id_mapper_io_req_valid),
    .io_req_ready(put_id_mapper_io_req_ready),
    .io_req_tl_id(put_id_mapper_io_req_tl_id),
    .io_req_nasti_id(put_id_mapper_io_req_nasti_id),
    .io_resp_valid(put_id_mapper_io_resp_valid),
    .io_resp_matches(put_id_mapper_io_resp_matches),
    .io_resp_nasti_id(put_id_mapper_io_resp_nasti_id),
    .io_resp_tl_id(put_id_mapper_io_resp_tl_id)
  );
  Arbiter_13 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_0_bits_client_id(gnt_arb_io_in_0_bits_client_id),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_1_bits_client_id(gnt_arb_io_in_1_bits_client_id),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_out_bits_client_id(gnt_arb_io_out_bits_client_id),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_tl_acquire_ready = T_955;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_nasti_aw_valid = T_865;
  assign io_nasti_aw_bits_addr = T_885_addr;
  assign io_nasti_aw_bits_len = T_885_len;
  assign io_nasti_aw_bits_size = T_885_size;
  assign io_nasti_aw_bits_burst = T_885_burst;
  assign io_nasti_aw_bits_lock = T_885_lock;
  assign io_nasti_aw_bits_cache = T_885_cache;
  assign io_nasti_aw_bits_prot = T_885_prot;
  assign io_nasti_aw_bits_qos = T_885_qos;
  assign io_nasti_aw_bits_region = T_885_region;
  assign io_nasti_aw_bits_id = T_885_id;
  assign io_nasti_aw_bits_user = T_885_user;
  assign io_nasti_w_valid = T_904;
  assign io_nasti_w_bits_data = T_940_data;
  assign io_nasti_w_bits_last = T_940_last;
  assign io_nasti_w_bits_id = T_940_id;
  assign io_nasti_w_bits_strb = T_940_strb;
  assign io_nasti_w_bits_user = T_940_user;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_ar_valid = T_789;
  assign io_nasti_ar_bits_addr = T_843_addr;
  assign io_nasti_ar_bits_len = T_843_len;
  assign io_nasti_ar_bits_size = T_843_size;
  assign io_nasti_ar_bits_burst = T_843_burst;
  assign io_nasti_ar_bits_lock = T_843_lock;
  assign io_nasti_ar_bits_cache = T_843_cache;
  assign io_nasti_ar_bits_prot = T_843_prot;
  assign io_nasti_ar_bits_qos = T_843_qos;
  assign io_nasti_ar_bits_region = T_843_region;
  assign io_nasti_ar_bits_id = T_843_id;
  assign io_nasti_ar_bits_user = T_843_user;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign T_688_0 = 3'h2;
  assign T_688_1 = 3'h3;
  assign T_688_2 = 3'h4;
  assign T_690 = T_688_0 == io_tl_acquire_bits_a_type;
  assign T_691 = T_688_1 == io_tl_acquire_bits_a_type;
  assign T_692 = T_688_2 == io_tl_acquire_bits_a_type;
  assign T_695 = T_690 | T_691;
  assign T_696 = T_695 | T_692;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T_696;
  assign T_705_0 = 3'h2;
  assign T_705_1 = 3'h0;
  assign T_705_2 = 3'h4;
  assign T_707 = T_705_0 == io_tl_acquire_bits_a_type;
  assign T_708 = T_705_1 == io_tl_acquire_bits_a_type;
  assign T_709 = T_705_2 == io_tl_acquire_bits_a_type;
  assign T_712 = T_707 | T_708;
  assign T_713 = T_712 | T_709;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T_713;
  assign T_722_0 = 3'h3;
  assign T_724 = T_722_0 == io_tl_acquire_bits_a_type;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T_724;
  assign T_727 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T_728 = T_727 & is_multibeat;
  assign T_731 = tl_cnt_out == 3'h7;
  assign GEN_6 = {{2'd0}, 1'h1};
  assign T_733 = tl_cnt_out + GEN_6;
  assign T_734 = T_733[2:0];
  assign GEN_0 = T_728 ? T_734 : tl_cnt_out;
  assign tl_wrap_out = T_728 & T_731;
  assign T_736 = has_data == 1'h0;
  assign get_valid = io_tl_acquire_valid & T_736;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign roq_clk = clk;
  assign roq_reset = reset;
  assign roq_io_enq_valid = T_776;
  assign roq_io_enq_bits_data_addr_beat = io_tl_acquire_bits_addr_beat;
  assign roq_io_enq_bits_data_subblock = is_subblock;
  assign roq_io_enq_bits_tag = io_nasti_ar_bits_id;
  assign roq_io_deq_valid = T_779;
  assign roq_io_deq_tag = io_nasti_r_bits_id;
  assign get_id_mapper_clk = clk;
  assign get_id_mapper_reset = reset;
  assign get_id_mapper_io_req_valid = T_781;
  assign get_id_mapper_io_req_tl_id = io_tl_acquire_bits_client_xact_id;
  assign get_id_mapper_io_resp_valid = T_783;
  assign get_id_mapper_io_resp_nasti_id = io_nasti_r_bits_id;
  assign put_id_mapper_clk = clk;
  assign put_id_mapper_reset = reset;
  assign put_id_mapper_io_req_valid = T_786;
  assign put_id_mapper_io_req_tl_id = io_tl_acquire_bits_client_xact_id;
  assign put_id_mapper_io_resp_valid = T_787;
  assign put_id_mapper_io_resp_nasti_id = io_nasti_b_bits_id;
  assign GEN_7 = {{2'd0}, 1'h0};
  assign T_761 = io_tl_acquire_bits_addr_beat == GEN_7;
  assign put_id_mask = is_subblock | T_761;
  assign T_763 = put_id_mask == 1'h0;
  assign put_id_ready = put_id_mapper_io_req_ready | T_763;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T_765 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_767 = roq_io_deq_data_subblock == 1'h0;
  assign T_768 = T_765 & T_767;
  assign T_771 = nasti_cnt_out == 3'h7;
  assign T_773 = nasti_cnt_out + GEN_6;
  assign T_774 = T_773[2:0];
  assign GEN_1 = T_768 ? T_774 : nasti_cnt_out;
  assign nasti_wrap_out = T_768 & T_771;
  assign T_775 = get_valid & io_nasti_ar_ready;
  assign T_776 = T_775 & get_id_mapper_io_req_ready;
  assign T_778 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign T_779 = T_765 & T_778;
  assign T_780 = get_valid & roq_io_enq_ready;
  assign T_781 = T_780 & io_nasti_ar_ready;
  assign T_783 = T_765 & io_nasti_r_bits_last;
  assign T_784 = put_valid & aw_ready;
  assign T_785 = T_784 & io_nasti_w_ready;
  assign T_786 = T_785 & put_id_mask;
  assign T_787 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_789 = T_780 & get_id_mapper_io_req_ready;
  assign T_790 = io_tl_acquire_bits_union[11:9];
  assign T_791 = {io_tl_acquire_bits_addr_block,io_tl_acquire_bits_addr_beat};
  assign T_792 = {T_791,T_790};
  assign T_793 = io_tl_acquire_bits_union[8:6];
  assign T_803 = 3'h7 == T_793;
  assign T_804 = T_803 ? {{1'd0}, 2'h3} : 3'h7;
  assign T_805 = 3'h3 == T_793;
  assign T_806 = T_805 ? {{1'd0}, 2'h3} : T_804;
  assign T_807 = 3'h6 == T_793;
  assign T_808 = T_807 ? {{1'd0}, 2'h2} : T_806;
  assign T_809 = 3'h2 == T_793;
  assign T_810 = T_809 ? {{1'd0}, 2'h2} : T_808;
  assign T_811 = 3'h5 == T_793;
  assign T_812 = T_811 ? {{2'd0}, 1'h1} : T_810;
  assign T_813 = 3'h1 == T_793;
  assign T_814 = T_813 ? {{2'd0}, 1'h1} : T_812;
  assign T_815 = 3'h4 == T_793;
  assign T_816 = T_815 ? {{2'd0}, 1'h0} : T_814;
  assign T_817 = 3'h0 == T_793;
  assign T_818 = T_817 ? {{2'd0}, 1'h0} : T_816;
  assign T_820 = is_subblock ? T_818 : {{1'd0}, 2'h3};
  assign T_823 = is_subblock ? {{2'd0}, 1'h0} : 3'h7;
  assign T_843_addr = T_792;
  assign T_843_len = {{5'd0}, T_823};
  assign T_843_size = T_820;
  assign T_843_burst = 2'h1;
  assign T_843_lock = 1'h0;
  assign T_843_cache = {{3'd0}, 1'h0};
  assign T_843_prot = {{2'd0}, 1'h0};
  assign T_843_qos = {{3'd0}, 1'h0};
  assign T_843_region = {{3'd0}, 1'h0};
  assign T_843_id = get_id_mapper_io_req_nasti_id;
  assign T_843_user = 1'h0;
  assign T_862 = w_inflight == 1'h0;
  assign T_863 = put_valid & io_nasti_w_ready;
  assign T_864 = T_863 & put_id_ready;
  assign T_865 = T_864 & T_862;
  assign T_872 = is_multibeat ? 3'h7 : {{2'd0}, 1'h0};
  assign T_885_addr = T_792;
  assign T_885_len = {{5'd0}, T_872};
  assign T_885_size = {{1'd0}, 2'h3};
  assign T_885_burst = 2'h1;
  assign T_885_lock = 1'h0;
  assign T_885_cache = 4'h0;
  assign T_885_prot = 3'h0;
  assign T_885_qos = 4'h0;
  assign T_885_region = 4'h0;
  assign T_885_id = put_id_mapper_io_req_nasti_id;
  assign T_885_user = 1'h0;
  assign T_904 = T_784 & put_id_ready;
  assign T_906 = io_tl_acquire_bits_a_type == 3'h4;
  assign T_907 = io_tl_acquire_bits_is_builtin_type & T_906;
  assign GEN_9 = {{7'd0}, 1'h1};
  assign T_911 = 8'h0 - GEN_9;
  assign T_912 = T_911[7:0];
  assign T_918_0 = T_912;
  assign T_921 = io_tl_acquire_bits_a_type == 3'h3;
  assign T_922 = io_tl_acquire_bits_is_builtin_type & T_921;
  assign T_924 = io_tl_acquire_bits_a_type == 3'h2;
  assign T_925 = io_tl_acquire_bits_is_builtin_type & T_924;
  assign T_926 = T_922 | T_925;
  assign T_927 = io_tl_acquire_bits_union[8:1];
  assign T_929 = T_926 ? T_927 : {{7'd0}, 1'h0};
  assign T_930 = T_907 ? T_918_0 : T_929;
  assign T_932 = T_727 & is_subblock;
  assign T_933 = tl_wrap_out | T_932;
  assign T_940_data = io_tl_acquire_bits_data;
  assign T_940_last = T_933;
  assign T_940_id = GEN_8;
  assign T_940_strb = T_930;
  assign T_940_user = 1'h0;
  assign T_951 = aw_ready & io_nasti_w_ready;
  assign T_952 = T_951 & put_id_ready;
  assign T_953 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T_954 = T_953 & get_id_mapper_io_req_ready;
  assign T_955 = has_data ? T_952 : T_954;
  assign T_959 = T_862 & T_727;
  assign T_960 = T_959 & is_multibeat;
  assign GEN_2 = T_960 ? 1'h1 : w_inflight;
  assign GEN_3 = tl_wrap_out ? 1'h0 : GEN_2;
  assign GEN_4 = w_inflight ? GEN_3 : GEN_2;
  assign T_963 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_971_0 = 3'h5;
  assign GEN_10 = {{1'd0}, T_971_0};
  assign T_973 = GEN_10 == io_tl_grant_bits_g_type;
  assign T_981_0 = 1'h0;
  assign GEN_11 = {{3'd0}, T_981_0};
  assign T_983 = GEN_11 == io_tl_grant_bits_g_type;
  assign T_986 = io_tl_grant_bits_is_builtin_type ? T_973 : T_983;
  assign T_988 = T_963 & T_986;
  assign T_993 = tl_cnt_in + GEN_6;
  assign T_994 = T_993[2:0];
  assign GEN_5 = T_988 ? T_994 : tl_cnt_in;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_nasti_r_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = T_1056_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = T_1056_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = T_1056_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = T_1056_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = T_1056_g_type;
  assign gnt_arb_io_in_0_bits_data = T_1056_data;
  assign gnt_arb_io_in_0_bits_client_id = GEN_12;
  assign gnt_arb_io_in_1_valid = io_nasti_b_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = T_1127_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = T_1127_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = T_1127_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = T_1127_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = T_1127_g_type;
  assign gnt_arb_io_in_1_bits_data = T_1127_data;
  assign gnt_arb_io_in_1_bits_client_id = GEN_14;
  assign gnt_arb_io_out_ready = io_tl_grant_ready;
  assign T_1026 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T_1028 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T_1056_addr_beat = T_1028;
  assign T_1056_client_xact_id = get_id_mapper_io_resp_tl_id;
  assign T_1056_manager_xact_id = 1'h0;
  assign T_1056_is_builtin_type = 1'h1;
  assign T_1056_g_type = {{1'd0}, T_1026};
  assign T_1056_data = io_nasti_r_bits_data;
  assign T_1084 = roq_io_deq_valid == 1'h0;
  assign T_1085 = T_1084 | roq_io_deq_matches;
  assign T_1086 = T_1085 | reset;
  assign T_1088 = T_1086 == 1'h0;
  assign T_1090 = gnt_arb_io_in_0_valid == 1'h0;
  assign T_1091 = T_1090 | get_id_mapper_io_resp_matches;
  assign T_1092 = T_1091 | reset;
  assign T_1094 = T_1092 == 1'h0;
  assign T_1127_addr_beat = {{2'd0}, 1'h0};
  assign T_1127_client_xact_id = put_id_mapper_io_resp_tl_id;
  assign T_1127_manager_xact_id = 1'h0;
  assign T_1127_is_builtin_type = 1'h1;
  assign T_1127_g_type = {{1'd0}, 3'h3};
  assign T_1127_data = {{63'd0}, 1'h0};
  assign T_1155 = gnt_arb_io_in_1_valid == 1'h0;
  assign T_1156 = T_1155 | put_id_mapper_io_resp_matches;
  assign T_1157 = T_1156 | reset;
  assign T_1159 = T_1157 == 1'h0;
  assign T_1161 = io_nasti_r_valid == 1'h0;
  assign GEN_13 = {{1'd0}, 1'h0};
  assign T_1163 = io_nasti_r_bits_resp == GEN_13;
  assign T_1164 = T_1161 | T_1163;
  assign T_1165 = T_1164 | reset;
  assign T_1167 = T_1165 == 1'h0;
  assign T_1169 = io_nasti_b_valid == 1'h0;
  assign T_1171 = io_nasti_b_bits_resp == GEN_13;
  assign T_1172 = T_1169 | T_1171;
  assign T_1173 = T_1172 | reset;
  assign T_1175 = T_1173 == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  tl_cnt_out = GEN_15[2:0];
  GEN_16 = {1{$random}};
  w_inflight = GEN_16[0:0];
  GEN_17 = {1{$random}};
  nasti_cnt_out = GEN_17[2:0];
  GEN_18 = {1{$random}};
  tl_cnt_in = GEN_18[2:0];
  GEN_19 = {1{$random}};
  GEN_8 = GEN_19[4:0];
  GEN_20 = {1{$random}};
  GEN_12 = GEN_20[0:0];
  GEN_21 = {1{$random}};
  GEN_14 = GEN_21[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else begin
      if(T_728) begin
        tl_cnt_out <= T_734;
      end
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else begin
      if(w_inflight) begin
        if(tl_wrap_out) begin
          w_inflight <= 1'h0;
        end else begin
          if(T_960) begin
            w_inflight <= 1'h1;
          end
        end
      end else begin
        if(T_960) begin
          w_inflight <= 1'h1;
        end
      end
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else begin
      if(T_768) begin
        nasti_cnt_out <= T_774;
      end
    end
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else begin
      if(T_988) begin
        tl_cnt_in <= T_994;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1088) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI converter ReorderQueue: NASTI tag error\n    at Nasti.scala:210 assert(!roq.io.deq.valid || roq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1088) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1088) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI ID Mapper: NASTI tag error\n    at Nasti.scala:212 assert(!gnt_arb.io.in(0).valid || get_id_mapper.io.resp.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1094) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1094) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1159) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at Nasti.scala:224 assert(!gnt_arb.io.in(1).valid || put_id_mapper.io.resp.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1159) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1167) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI read error\n    at Nasti.scala:226 assert(!io.nasti.r.valid || io.nasti.r.bits.resp === UInt(0), \"NASTI read error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1167) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1175) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI write error\n    at Nasti.scala:227 assert(!io.nasti.b.valid || io.nasti.b.bits.resp === UInt(0), \"NASTI write error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1175) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_15(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0] io_enq_bits_len,
  input  [2:0] io_enq_bits_size,
  input  [1:0] io_enq_bits_burst,
  input   io_enq_bits_lock,
  input  [3:0] io_enq_bits_cache,
  input  [2:0] io_enq_bits_prot,
  input  [3:0] io_enq_bits_qos,
  input  [3:0] io_enq_bits_region,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst,
  output  io_deq_bits_lock,
  output [3:0] io_deq_bits_cache,
  output [2:0] io_deq_bits_prot,
  output [3:0] io_deq_bits_qos,
  output [3:0] io_deq_bits_region,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [31:0] ram_addr [0:0];
  reg [31:0] GEN_0;
  wire [31:0] ram_addr_T_144_data;
  wire  ram_addr_T_144_addr;
  wire  ram_addr_T_144_en;
  wire [31:0] ram_addr_T_125_data;
  wire  ram_addr_T_125_addr;
  wire  ram_addr_T_125_mask;
  wire  ram_addr_T_125_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] GEN_1;
  wire [7:0] ram_len_T_144_data;
  wire  ram_len_T_144_addr;
  wire  ram_len_T_144_en;
  wire [7:0] ram_len_T_125_data;
  wire  ram_len_T_125_addr;
  wire  ram_len_T_125_mask;
  wire  ram_len_T_125_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_size_T_144_data;
  wire  ram_size_T_144_addr;
  wire  ram_size_T_144_en;
  wire [2:0] ram_size_T_125_data;
  wire  ram_size_T_125_addr;
  wire  ram_size_T_125_mask;
  wire  ram_size_T_125_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_burst_T_144_data;
  wire  ram_burst_T_144_addr;
  wire  ram_burst_T_144_en;
  wire [1:0] ram_burst_T_125_data;
  wire  ram_burst_T_125_addr;
  wire  ram_burst_T_125_mask;
  wire  ram_burst_T_125_en;
  reg  ram_lock [0:0];
  reg [31:0] GEN_4;
  wire  ram_lock_T_144_data;
  wire  ram_lock_T_144_addr;
  wire  ram_lock_T_144_en;
  wire  ram_lock_T_125_data;
  wire  ram_lock_T_125_addr;
  wire  ram_lock_T_125_mask;
  wire  ram_lock_T_125_en;
  reg [3:0] ram_cache [0:0];
  reg [31:0] GEN_5;
  wire [3:0] ram_cache_T_144_data;
  wire  ram_cache_T_144_addr;
  wire  ram_cache_T_144_en;
  wire [3:0] ram_cache_T_125_data;
  wire  ram_cache_T_125_addr;
  wire  ram_cache_T_125_mask;
  wire  ram_cache_T_125_en;
  reg [2:0] ram_prot [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_prot_T_144_data;
  wire  ram_prot_T_144_addr;
  wire  ram_prot_T_144_en;
  wire [2:0] ram_prot_T_125_data;
  wire  ram_prot_T_125_addr;
  wire  ram_prot_T_125_mask;
  wire  ram_prot_T_125_en;
  reg [3:0] ram_qos [0:0];
  reg [31:0] GEN_7;
  wire [3:0] ram_qos_T_144_data;
  wire  ram_qos_T_144_addr;
  wire  ram_qos_T_144_en;
  wire [3:0] ram_qos_T_125_data;
  wire  ram_qos_T_125_addr;
  wire  ram_qos_T_125_mask;
  wire  ram_qos_T_125_en;
  reg [3:0] ram_region [0:0];
  reg [31:0] GEN_8;
  wire [3:0] ram_region_T_144_data;
  wire  ram_region_T_144_addr;
  wire  ram_region_T_144_en;
  wire [3:0] ram_region_T_125_data;
  wire  ram_region_T_125_addr;
  wire  ram_region_T_125_mask;
  wire  ram_region_T_125_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_9;
  wire [4:0] ram_id_T_144_data;
  wire  ram_id_T_144_addr;
  wire  ram_id_T_144_en;
  wire [4:0] ram_id_T_125_data;
  wire  ram_id_T_125_addr;
  wire  ram_id_T_125_mask;
  wire  ram_id_T_125_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_10;
  wire  ram_user_T_144_data;
  wire  ram_user_T_144_addr;
  wire  ram_user_T_144_en;
  wire  ram_user_T_125_data;
  wire  ram_user_T_125_addr;
  wire  ram_user_T_125_mask;
  wire  ram_user_T_125_en;
  reg  maybe_full;
  reg [31:0] GEN_11;
  wire  T_122;
  wire  T_123;
  wire  do_enq;
  wire  T_124;
  wire  do_deq;
  wire  T_139;
  wire  GEN_25;
  wire  T_141;
  wire [1:0] T_156;
  wire  ptr_diff;
  wire [1:0] T_158;
  assign io_enq_ready = T_122;
  assign io_deq_valid = T_141;
  assign io_deq_bits_addr = ram_addr_T_144_data;
  assign io_deq_bits_len = ram_len_T_144_data;
  assign io_deq_bits_size = ram_size_T_144_data;
  assign io_deq_bits_burst = ram_burst_T_144_data;
  assign io_deq_bits_lock = ram_lock_T_144_data;
  assign io_deq_bits_cache = ram_cache_T_144_data;
  assign io_deq_bits_prot = ram_prot_T_144_data;
  assign io_deq_bits_qos = ram_qos_T_144_data;
  assign io_deq_bits_region = ram_region_T_144_data;
  assign io_deq_bits_id = ram_id_T_144_data;
  assign io_deq_bits_user = ram_user_T_144_data;
  assign io_count = T_158[0];
  assign ram_addr_T_144_addr = 1'h0;
  assign ram_addr_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_T_144_data = ram_addr[ram_addr_T_144_addr];
  `else
  assign ram_addr_T_144_data = ram_addr_T_144_addr >= 1'h1 ? $random : ram_addr[ram_addr_T_144_addr];
  `endif
  assign ram_addr_T_125_data = io_enq_bits_addr;
  assign ram_addr_T_125_addr = 1'h0;
  assign ram_addr_T_125_mask = do_enq;
  assign ram_addr_T_125_en = do_enq;
  assign ram_len_T_144_addr = 1'h0;
  assign ram_len_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_len_T_144_data = ram_len[ram_len_T_144_addr];
  `else
  assign ram_len_T_144_data = ram_len_T_144_addr >= 1'h1 ? $random : ram_len[ram_len_T_144_addr];
  `endif
  assign ram_len_T_125_data = io_enq_bits_len;
  assign ram_len_T_125_addr = 1'h0;
  assign ram_len_T_125_mask = do_enq;
  assign ram_len_T_125_en = do_enq;
  assign ram_size_T_144_addr = 1'h0;
  assign ram_size_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_size_T_144_data = ram_size[ram_size_T_144_addr];
  `else
  assign ram_size_T_144_data = ram_size_T_144_addr >= 1'h1 ? $random : ram_size[ram_size_T_144_addr];
  `endif
  assign ram_size_T_125_data = io_enq_bits_size;
  assign ram_size_T_125_addr = 1'h0;
  assign ram_size_T_125_mask = do_enq;
  assign ram_size_T_125_en = do_enq;
  assign ram_burst_T_144_addr = 1'h0;
  assign ram_burst_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_burst_T_144_data = ram_burst[ram_burst_T_144_addr];
  `else
  assign ram_burst_T_144_data = ram_burst_T_144_addr >= 1'h1 ? $random : ram_burst[ram_burst_T_144_addr];
  `endif
  assign ram_burst_T_125_data = io_enq_bits_burst;
  assign ram_burst_T_125_addr = 1'h0;
  assign ram_burst_T_125_mask = do_enq;
  assign ram_burst_T_125_en = do_enq;
  assign ram_lock_T_144_addr = 1'h0;
  assign ram_lock_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_lock_T_144_data = ram_lock[ram_lock_T_144_addr];
  `else
  assign ram_lock_T_144_data = ram_lock_T_144_addr >= 1'h1 ? $random : ram_lock[ram_lock_T_144_addr];
  `endif
  assign ram_lock_T_125_data = io_enq_bits_lock;
  assign ram_lock_T_125_addr = 1'h0;
  assign ram_lock_T_125_mask = do_enq;
  assign ram_lock_T_125_en = do_enq;
  assign ram_cache_T_144_addr = 1'h0;
  assign ram_cache_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_cache_T_144_data = ram_cache[ram_cache_T_144_addr];
  `else
  assign ram_cache_T_144_data = ram_cache_T_144_addr >= 1'h1 ? $random : ram_cache[ram_cache_T_144_addr];
  `endif
  assign ram_cache_T_125_data = io_enq_bits_cache;
  assign ram_cache_T_125_addr = 1'h0;
  assign ram_cache_T_125_mask = do_enq;
  assign ram_cache_T_125_en = do_enq;
  assign ram_prot_T_144_addr = 1'h0;
  assign ram_prot_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_prot_T_144_data = ram_prot[ram_prot_T_144_addr];
  `else
  assign ram_prot_T_144_data = ram_prot_T_144_addr >= 1'h1 ? $random : ram_prot[ram_prot_T_144_addr];
  `endif
  assign ram_prot_T_125_data = io_enq_bits_prot;
  assign ram_prot_T_125_addr = 1'h0;
  assign ram_prot_T_125_mask = do_enq;
  assign ram_prot_T_125_en = do_enq;
  assign ram_qos_T_144_addr = 1'h0;
  assign ram_qos_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_qos_T_144_data = ram_qos[ram_qos_T_144_addr];
  `else
  assign ram_qos_T_144_data = ram_qos_T_144_addr >= 1'h1 ? $random : ram_qos[ram_qos_T_144_addr];
  `endif
  assign ram_qos_T_125_data = io_enq_bits_qos;
  assign ram_qos_T_125_addr = 1'h0;
  assign ram_qos_T_125_mask = do_enq;
  assign ram_qos_T_125_en = do_enq;
  assign ram_region_T_144_addr = 1'h0;
  assign ram_region_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_region_T_144_data = ram_region[ram_region_T_144_addr];
  `else
  assign ram_region_T_144_data = ram_region_T_144_addr >= 1'h1 ? $random : ram_region[ram_region_T_144_addr];
  `endif
  assign ram_region_T_125_data = io_enq_bits_region;
  assign ram_region_T_125_addr = 1'h0;
  assign ram_region_T_125_mask = do_enq;
  assign ram_region_T_125_en = do_enq;
  assign ram_id_T_144_addr = 1'h0;
  assign ram_id_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_id_T_144_data = ram_id[ram_id_T_144_addr];
  `else
  assign ram_id_T_144_data = ram_id_T_144_addr >= 1'h1 ? $random : ram_id[ram_id_T_144_addr];
  `endif
  assign ram_id_T_125_data = io_enq_bits_id;
  assign ram_id_T_125_addr = 1'h0;
  assign ram_id_T_125_mask = do_enq;
  assign ram_id_T_125_en = do_enq;
  assign ram_user_T_144_addr = 1'h0;
  assign ram_user_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_user_T_144_data = ram_user[ram_user_T_144_addr];
  `else
  assign ram_user_T_144_data = ram_user_T_144_addr >= 1'h1 ? $random : ram_user[ram_user_T_144_addr];
  `endif
  assign ram_user_T_125_data = io_enq_bits_user;
  assign ram_user_T_125_addr = 1'h0;
  assign ram_user_T_125_mask = do_enq;
  assign ram_user_T_125_en = do_enq;
  assign T_122 = maybe_full == 1'h0;
  assign T_123 = io_enq_ready & io_enq_valid;
  assign do_enq = T_123;
  assign T_124 = io_deq_ready & io_deq_valid;
  assign do_deq = T_124;
  assign T_139 = do_enq != do_deq;
  assign GEN_25 = T_139 ? do_enq : maybe_full;
  assign T_141 = T_122 == 1'h0;
  assign T_156 = 1'h0 - 1'h0;
  assign ptr_diff = T_156[0:0];
  assign T_158 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = GEN_0[31:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = GEN_1[7:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = GEN_2[2:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = GEN_3[1:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_lock[initvar] = GEN_4[0:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = GEN_5[3:0];
  GEN_6 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = GEN_6[2:0];
  GEN_7 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_qos[initvar] = GEN_7[3:0];
  GEN_8 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_region[initvar] = GEN_8[3:0];
  GEN_9 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_9[4:0];
  GEN_10 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_10[0:0];
  GEN_11 = {1{$random}};
  maybe_full = GEN_11[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_T_125_en & ram_addr_T_125_mask) begin
      ram_addr[ram_addr_T_125_addr] <= ram_addr_T_125_data;
    end
    if(ram_len_T_125_en & ram_len_T_125_mask) begin
      ram_len[ram_len_T_125_addr] <= ram_len_T_125_data;
    end
    if(ram_size_T_125_en & ram_size_T_125_mask) begin
      ram_size[ram_size_T_125_addr] <= ram_size_T_125_data;
    end
    if(ram_burst_T_125_en & ram_burst_T_125_mask) begin
      ram_burst[ram_burst_T_125_addr] <= ram_burst_T_125_data;
    end
    if(ram_lock_T_125_en & ram_lock_T_125_mask) begin
      ram_lock[ram_lock_T_125_addr] <= ram_lock_T_125_data;
    end
    if(ram_cache_T_125_en & ram_cache_T_125_mask) begin
      ram_cache[ram_cache_T_125_addr] <= ram_cache_T_125_data;
    end
    if(ram_prot_T_125_en & ram_prot_T_125_mask) begin
      ram_prot[ram_prot_T_125_addr] <= ram_prot_T_125_data;
    end
    if(ram_qos_T_125_en & ram_qos_T_125_mask) begin
      ram_qos[ram_qos_T_125_addr] <= ram_qos_T_125_data;
    end
    if(ram_region_T_125_en & ram_region_T_125_mask) begin
      ram_region[ram_region_T_125_addr] <= ram_region_T_125_data;
    end
    if(ram_id_T_125_en & ram_id_T_125_mask) begin
      ram_id[ram_id_T_125_addr] <= ram_id_T_125_data;
    end
    if(ram_user_T_125_en & ram_user_T_125_mask) begin
      ram_user[ram_user_T_125_addr] <= ram_user_T_125_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_17(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input  [7:0] io_enq_bits_strb,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output [7:0] io_deq_bits_strb,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_0;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_1;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_2;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg [7:0] ram_strb [0:1];
  reg [31:0] GEN_3;
  wire [7:0] ram_strb_T_94_data;
  wire  ram_strb_T_94_addr;
  wire  ram_strb_T_94_en;
  wire [7:0] ram_strb_T_73_data;
  wire  ram_strb_T_73_addr;
  wire  ram_strb_T_73_mask;
  wire  ram_strb_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_strb = ram_strb_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  `else
  assign ram_data_T_94_data = ram_data_T_94_addr >= 2'h2 ? $random : ram_data[ram_data_T_94_addr];
  `endif
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  `else
  assign ram_last_T_94_data = ram_last_T_94_addr >= 2'h2 ? $random : ram_last[ram_last_T_94_addr];
  `endif
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  `else
  assign ram_id_T_94_data = ram_id_T_94_addr >= 2'h2 ? $random : ram_id[ram_id_T_94_addr];
  `endif
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_strb_T_94_addr = T_67;
  assign ram_strb_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_strb_T_94_data = ram_strb[ram_strb_T_94_addr];
  `else
  assign ram_strb_T_94_data = ram_strb_T_94_addr >= 2'h2 ? $random : ram_strb[ram_strb_T_94_addr];
  `endif
  assign ram_strb_T_73_data = io_enq_bits_strb;
  assign ram_strb_T_73_addr = T_65;
  assign ram_strb_T_73_mask = do_enq;
  assign ram_strb_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  `else
  assign ram_user_T_94_data = ram_user_T_94_addr >= 2'h2 ? $random : ram_user[ram_user_T_94_addr];
  `endif
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {2{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_0[63:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_1[0:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_2[4:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = GEN_3[7:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_strb_T_73_en & ram_strb_T_73_mask) begin
      ram_strb[ram_strb_T_73_addr] <= ram_strb_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_65 <= T_83;
      end
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_67 <= T_88;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_89) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_18(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [1:0] ram_resp [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_94_data;
  wire  ram_resp_T_94_addr;
  wire  ram_resp_T_94_en;
  wire [1:0] ram_resp_T_73_data;
  wire  ram_resp_T_73_addr;
  wire  ram_resp_T_73_mask;
  wire  ram_resp_T_73_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_1;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_2;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_3;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_resp = ram_resp_T_94_data;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_resp_T_94_addr = T_67;
  assign ram_resp_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_resp_T_94_data = ram_resp[ram_resp_T_94_addr];
  `else
  assign ram_resp_T_94_data = ram_resp_T_94_addr >= 2'h2 ? $random : ram_resp[ram_resp_T_94_addr];
  `endif
  assign ram_resp_T_73_data = io_enq_bits_resp;
  assign ram_resp_T_73_addr = T_65;
  assign ram_resp_T_73_mask = do_enq;
  assign ram_resp_T_73_en = do_enq;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  `else
  assign ram_data_T_94_data = ram_data_T_94_addr >= 2'h2 ? $random : ram_data[ram_data_T_94_addr];
  `endif
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  `else
  assign ram_last_T_94_data = ram_last_T_94_addr >= 2'h2 ? $random : ram_last[ram_last_T_94_addr];
  `endif
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  `else
  assign ram_id_T_94_data = ram_id_T_94_addr >= 2'h2 ? $random : ram_id[ram_id_T_94_addr];
  `endif
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  `else
  assign ram_user_T_94_data = ram_user_T_94_addr >= 2'h2 ? $random : ram_user[ram_user_T_94_addr];
  `endif
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  GEN_1 = {2{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_1[63:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_2[0:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_3[4:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_73_en & ram_resp_T_73_mask) begin
      ram_resp[ram_resp_T_73_addr] <= ram_resp_T_73_data;
    end
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_65 <= T_83;
      end
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_67 <= T_88;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_89) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_19(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [1:0] ram_resp [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_64_data;
  wire  ram_resp_T_64_addr;
  wire  ram_resp_T_64_en;
  wire [1:0] ram_resp_T_53_data;
  wire  ram_resp_T_53_addr;
  wire  ram_resp_T_53_mask;
  wire  ram_resp_T_53_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_1;
  wire [4:0] ram_id_T_64_data;
  wire  ram_id_T_64_addr;
  wire  ram_id_T_64_en;
  wire [4:0] ram_id_T_53_data;
  wire  ram_id_T_53_addr;
  wire  ram_id_T_53_mask;
  wire  ram_id_T_53_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_2;
  wire  ram_user_T_64_data;
  wire  ram_user_T_64_addr;
  wire  ram_user_T_64_en;
  wire  ram_user_T_53_data;
  wire  ram_user_T_53_addr;
  wire  ram_user_T_53_mask;
  wire  ram_user_T_53_en;
  reg  maybe_full;
  reg [31:0] GEN_3;
  wire  T_50;
  wire  T_51;
  wire  do_enq;
  wire  T_52;
  wire  do_deq;
  wire  T_59;
  wire  GEN_9;
  wire  T_61;
  wire [1:0] T_68;
  wire  ptr_diff;
  wire [1:0] T_70;
  assign io_enq_ready = T_50;
  assign io_deq_valid = T_61;
  assign io_deq_bits_resp = ram_resp_T_64_data;
  assign io_deq_bits_id = ram_id_T_64_data;
  assign io_deq_bits_user = ram_user_T_64_data;
  assign io_count = T_70[0];
  assign ram_resp_T_64_addr = 1'h0;
  assign ram_resp_T_64_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_resp_T_64_data = ram_resp[ram_resp_T_64_addr];
  `else
  assign ram_resp_T_64_data = ram_resp_T_64_addr >= 1'h1 ? $random : ram_resp[ram_resp_T_64_addr];
  `endif
  assign ram_resp_T_53_data = io_enq_bits_resp;
  assign ram_resp_T_53_addr = 1'h0;
  assign ram_resp_T_53_mask = do_enq;
  assign ram_resp_T_53_en = do_enq;
  assign ram_id_T_64_addr = 1'h0;
  assign ram_id_T_64_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_id_T_64_data = ram_id[ram_id_T_64_addr];
  `else
  assign ram_id_T_64_data = ram_id_T_64_addr >= 1'h1 ? $random : ram_id[ram_id_T_64_addr];
  `endif
  assign ram_id_T_53_data = io_enq_bits_id;
  assign ram_id_T_53_addr = 1'h0;
  assign ram_id_T_53_mask = do_enq;
  assign ram_id_T_53_en = do_enq;
  assign ram_user_T_64_addr = 1'h0;
  assign ram_user_T_64_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_user_T_64_data = ram_user[ram_user_T_64_addr];
  `else
  assign ram_user_T_64_data = ram_user_T_64_addr >= 1'h1 ? $random : ram_user[ram_user_T_64_addr];
  `endif
  assign ram_user_T_53_data = io_enq_bits_user;
  assign ram_user_T_53_addr = 1'h0;
  assign ram_user_T_53_mask = do_enq;
  assign ram_user_T_53_en = do_enq;
  assign T_50 = maybe_full == 1'h0;
  assign T_51 = io_enq_ready & io_enq_valid;
  assign do_enq = T_51;
  assign T_52 = io_deq_ready & io_deq_valid;
  assign do_deq = T_52;
  assign T_59 = do_enq != do_deq;
  assign GEN_9 = T_59 ? do_enq : maybe_full;
  assign T_61 = T_50 == 1'h0;
  assign T_68 = 1'h0 - 1'h0;
  assign ptr_diff = T_68[0:0];
  assign T_70 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_1[4:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_2[0:0];
  GEN_3 = {1{$random}};
  maybe_full = GEN_3[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_53_en & ram_resp_T_53_mask) begin
      ram_resp[ram_resp_T_53_addr] <= ram_resp_T_53_data;
    end
    if(ram_id_T_53_en & ram_id_T_53_mask) begin
      ram_id[ram_id_T_53_addr] <= ram_id_T_53_data;
    end
    if(ram_user_T_53_en & ram_user_T_53_mask) begin
      ram_user[ram_user_T_53_addr] <= ram_user_T_53_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_59) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module OuterMemorySystem(
  input   clk,
  input   reset,
  output  io_tiles_cached_0_acquire_ready,
  input   io_tiles_cached_0_acquire_valid,
  input  [25:0] io_tiles_cached_0_acquire_bits_addr_block,
  input  [1:0] io_tiles_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_cached_0_acquire_bits_addr_beat,
  input   io_tiles_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_cached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_cached_0_acquire_bits_union,
  input  [63:0] io_tiles_cached_0_acquire_bits_data,
  input   io_tiles_cached_0_probe_ready,
  output  io_tiles_cached_0_probe_valid,
  output [25:0] io_tiles_cached_0_probe_bits_addr_block,
  output [1:0] io_tiles_cached_0_probe_bits_p_type,
  output  io_tiles_cached_0_release_ready,
  input   io_tiles_cached_0_release_valid,
  input  [2:0] io_tiles_cached_0_release_bits_addr_beat,
  input  [25:0] io_tiles_cached_0_release_bits_addr_block,
  input  [1:0] io_tiles_cached_0_release_bits_client_xact_id,
  input   io_tiles_cached_0_release_bits_voluntary,
  input  [2:0] io_tiles_cached_0_release_bits_r_type,
  input  [63:0] io_tiles_cached_0_release_bits_data,
  input   io_tiles_cached_0_grant_ready,
  output  io_tiles_cached_0_grant_valid,
  output [2:0] io_tiles_cached_0_grant_bits_addr_beat,
  output [1:0] io_tiles_cached_0_grant_bits_client_xact_id,
  output [2:0] io_tiles_cached_0_grant_bits_manager_xact_id,
  output  io_tiles_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_cached_0_grant_bits_g_type,
  output [63:0] io_tiles_cached_0_grant_bits_data,
  output  io_tiles_cached_0_grant_bits_manager_id,
  output  io_tiles_cached_0_finish_ready,
  input   io_tiles_cached_0_finish_valid,
  input  [2:0] io_tiles_cached_0_finish_bits_manager_xact_id,
  input   io_tiles_cached_0_finish_bits_manager_id,
  output  io_tiles_uncached_0_acquire_ready,
  input   io_tiles_uncached_0_acquire_valid,
  input  [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
  input  [1:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_uncached_0_acquire_bits_addr_beat,
  input   io_tiles_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_uncached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_uncached_0_acquire_bits_union,
  input  [63:0] io_tiles_uncached_0_acquire_bits_data,
  input   io_tiles_uncached_0_grant_ready,
  output  io_tiles_uncached_0_grant_valid,
  output [2:0] io_tiles_uncached_0_grant_bits_addr_beat,
  output [1:0] io_tiles_uncached_0_grant_bits_client_xact_id,
  output [2:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
  output  io_tiles_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_uncached_0_grant_bits_g_type,
  output [63:0] io_tiles_uncached_0_grant_bits_data,
  input   io_incoherent_0,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  input   io_mmio_acquire_ready,
  output  io_mmio_acquire_valid,
  output [25:0] io_mmio_acquire_bits_addr_block,
  output [1:0] io_mmio_acquire_bits_client_xact_id,
  output [2:0] io_mmio_acquire_bits_addr_beat,
  output  io_mmio_acquire_bits_is_builtin_type,
  output [2:0] io_mmio_acquire_bits_a_type,
  output [11:0] io_mmio_acquire_bits_union,
  output [63:0] io_mmio_acquire_bits_data,
  output  io_mmio_grant_ready,
  input   io_mmio_grant_valid,
  input  [2:0] io_mmio_grant_bits_addr_beat,
  input  [1:0] io_mmio_grant_bits_client_xact_id,
  input   io_mmio_grant_bits_manager_xact_id,
  input   io_mmio_grant_bits_is_builtin_type,
  input  [3:0] io_mmio_grant_bits_g_type,
  input  [63:0] io_mmio_grant_bits_data
);
  wire  l1tol2net_clk;
  wire  l1tol2net_reset;
  wire  l1tol2net_io_clients_cached_0_acquire_ready;
  wire  l1tol2net_io_clients_cached_0_acquire_valid;
  wire [25:0] l1tol2net_io_clients_cached_0_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_cached_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_clients_cached_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_clients_cached_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_clients_cached_0_acquire_bits_data;
  wire  l1tol2net_io_clients_cached_0_probe_ready;
  wire  l1tol2net_io_clients_cached_0_probe_valid;
  wire [25:0] l1tol2net_io_clients_cached_0_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_cached_0_probe_bits_p_type;
  wire  l1tol2net_io_clients_cached_0_release_ready;
  wire  l1tol2net_io_clients_cached_0_release_valid;
  wire [2:0] l1tol2net_io_clients_cached_0_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_clients_cached_0_release_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_cached_0_release_bits_client_xact_id;
  wire  l1tol2net_io_clients_cached_0_release_bits_voluntary;
  wire [2:0] l1tol2net_io_clients_cached_0_release_bits_r_type;
  wire [63:0] l1tol2net_io_clients_cached_0_release_bits_data;
  wire  l1tol2net_io_clients_cached_0_grant_ready;
  wire  l1tol2net_io_clients_cached_0_grant_valid;
  wire [2:0] l1tol2net_io_clients_cached_0_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_clients_cached_0_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_clients_cached_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_clients_cached_0_grant_bits_data;
  wire  l1tol2net_io_clients_cached_0_grant_bits_manager_id;
  wire  l1tol2net_io_clients_cached_0_finish_ready;
  wire  l1tol2net_io_clients_cached_0_finish_valid;
  wire [2:0] l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id;
  wire  l1tol2net_io_clients_cached_0_finish_bits_manager_id;
  wire  l1tol2net_io_clients_uncached_0_acquire_ready;
  wire  l1tol2net_io_clients_uncached_0_acquire_valid;
  wire [25:0] l1tol2net_io_clients_uncached_0_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_clients_uncached_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_clients_uncached_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_clients_uncached_0_acquire_bits_data;
  wire  l1tol2net_io_clients_uncached_0_grant_ready;
  wire  l1tol2net_io_clients_uncached_0_grant_valid;
  wire [2:0] l1tol2net_io_clients_uncached_0_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_clients_uncached_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_clients_uncached_0_grant_bits_data;
  wire  l1tol2net_io_managers_0_acquire_ready;
  wire  l1tol2net_io_managers_0_acquire_valid;
  wire [25:0] l1tol2net_io_managers_0_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_managers_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_managers_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_managers_0_acquire_bits_data;
  wire  l1tol2net_io_managers_0_acquire_bits_client_id;
  wire  l1tol2net_io_managers_0_grant_ready;
  wire  l1tol2net_io_managers_0_grant_valid;
  wire [2:0] l1tol2net_io_managers_0_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_managers_0_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_managers_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_managers_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_managers_0_grant_bits_data;
  wire  l1tol2net_io_managers_0_grant_bits_client_id;
  wire  l1tol2net_io_managers_0_finish_ready;
  wire  l1tol2net_io_managers_0_finish_valid;
  wire [2:0] l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  wire  l1tol2net_io_managers_0_probe_ready;
  wire  l1tol2net_io_managers_0_probe_valid;
  wire [25:0] l1tol2net_io_managers_0_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_0_probe_bits_p_type;
  wire  l1tol2net_io_managers_0_probe_bits_client_id;
  wire  l1tol2net_io_managers_0_release_ready;
  wire  l1tol2net_io_managers_0_release_valid;
  wire [2:0] l1tol2net_io_managers_0_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_managers_0_release_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_0_release_bits_client_xact_id;
  wire  l1tol2net_io_managers_0_release_bits_voluntary;
  wire [2:0] l1tol2net_io_managers_0_release_bits_r_type;
  wire [63:0] l1tol2net_io_managers_0_release_bits_data;
  wire  l1tol2net_io_managers_0_release_bits_client_id;
  wire  l1tol2net_io_managers_1_acquire_ready;
  wire  l1tol2net_io_managers_1_acquire_valid;
  wire [25:0] l1tol2net_io_managers_1_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_1_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_1_acquire_bits_addr_beat;
  wire  l1tol2net_io_managers_1_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_managers_1_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_managers_1_acquire_bits_union;
  wire [63:0] l1tol2net_io_managers_1_acquire_bits_data;
  wire  l1tol2net_io_managers_1_acquire_bits_client_id;
  wire  l1tol2net_io_managers_1_grant_ready;
  wire  l1tol2net_io_managers_1_grant_valid;
  wire [2:0] l1tol2net_io_managers_1_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_managers_1_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_1_grant_bits_manager_xact_id;
  wire  l1tol2net_io_managers_1_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_managers_1_grant_bits_g_type;
  wire [63:0] l1tol2net_io_managers_1_grant_bits_data;
  wire  l1tol2net_io_managers_1_grant_bits_client_id;
  wire  l1tol2net_io_managers_1_finish_ready;
  wire  l1tol2net_io_managers_1_finish_valid;
  wire [2:0] l1tol2net_io_managers_1_finish_bits_manager_xact_id;
  wire  l1tol2net_io_managers_1_probe_ready;
  wire  l1tol2net_io_managers_1_probe_valid;
  wire [25:0] l1tol2net_io_managers_1_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_1_probe_bits_p_type;
  wire  l1tol2net_io_managers_1_probe_bits_client_id;
  wire  l1tol2net_io_managers_1_release_ready;
  wire  l1tol2net_io_managers_1_release_valid;
  wire [2:0] l1tol2net_io_managers_1_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_managers_1_release_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_1_release_bits_client_xact_id;
  wire  l1tol2net_io_managers_1_release_bits_voluntary;
  wire [2:0] l1tol2net_io_managers_1_release_bits_r_type;
  wire [63:0] l1tol2net_io_managers_1_release_bits_data;
  wire  l1tol2net_io_managers_1_release_bits_client_id;
  wire  L2BroadcastHub_1_clk;
  wire  L2BroadcastHub_1_reset;
  wire  L2BroadcastHub_1_io_inner_acquire_ready;
  wire  L2BroadcastHub_1_io_inner_acquire_valid;
  wire [25:0] L2BroadcastHub_1_io_inner_acquire_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_1_io_inner_acquire_bits_addr_beat;
  wire  L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] L2BroadcastHub_1_io_inner_acquire_bits_a_type;
  wire [11:0] L2BroadcastHub_1_io_inner_acquire_bits_union;
  wire [63:0] L2BroadcastHub_1_io_inner_acquire_bits_data;
  wire  L2BroadcastHub_1_io_inner_acquire_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_grant_ready;
  wire  L2BroadcastHub_1_io_inner_grant_valid;
  wire [2:0] L2BroadcastHub_1_io_inner_grant_bits_addr_beat;
  wire [1:0] L2BroadcastHub_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] L2BroadcastHub_1_io_inner_grant_bits_g_type;
  wire [63:0] L2BroadcastHub_1_io_inner_grant_bits_data;
  wire  L2BroadcastHub_1_io_inner_grant_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_finish_ready;
  wire  L2BroadcastHub_1_io_inner_finish_valid;
  wire [2:0] L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_inner_probe_ready;
  wire  L2BroadcastHub_1_io_inner_probe_valid;
  wire [25:0] L2BroadcastHub_1_io_inner_probe_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_inner_probe_bits_p_type;
  wire  L2BroadcastHub_1_io_inner_probe_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_release_ready;
  wire  L2BroadcastHub_1_io_inner_release_valid;
  wire [2:0] L2BroadcastHub_1_io_inner_release_bits_addr_beat;
  wire [25:0] L2BroadcastHub_1_io_inner_release_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_inner_release_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_inner_release_bits_voluntary;
  wire [2:0] L2BroadcastHub_1_io_inner_release_bits_r_type;
  wire [63:0] L2BroadcastHub_1_io_inner_release_bits_data;
  wire  L2BroadcastHub_1_io_inner_release_bits_client_id;
  wire  L2BroadcastHub_1_io_incoherent_0;
  wire  L2BroadcastHub_1_io_outer_acquire_ready;
  wire  L2BroadcastHub_1_io_outer_acquire_valid;
  wire [25:0] L2BroadcastHub_1_io_outer_acquire_bits_addr_block;
  wire [2:0] L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_1_io_outer_acquire_bits_addr_beat;
  wire  L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] L2BroadcastHub_1_io_outer_acquire_bits_a_type;
  wire [11:0] L2BroadcastHub_1_io_outer_acquire_bits_union;
  wire [63:0] L2BroadcastHub_1_io_outer_acquire_bits_data;
  wire  L2BroadcastHub_1_io_outer_probe_ready;
  wire  L2BroadcastHub_1_io_outer_probe_valid;
  wire [25:0] L2BroadcastHub_1_io_outer_probe_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_outer_probe_bits_p_type;
  wire  L2BroadcastHub_1_io_outer_release_ready;
  wire  L2BroadcastHub_1_io_outer_release_valid;
  wire [2:0] L2BroadcastHub_1_io_outer_release_bits_addr_beat;
  wire [25:0] L2BroadcastHub_1_io_outer_release_bits_addr_block;
  wire [2:0] L2BroadcastHub_1_io_outer_release_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_outer_release_bits_voluntary;
  wire [2:0] L2BroadcastHub_1_io_outer_release_bits_r_type;
  wire [63:0] L2BroadcastHub_1_io_outer_release_bits_data;
  wire  L2BroadcastHub_1_io_outer_grant_ready;
  wire  L2BroadcastHub_1_io_outer_grant_valid;
  wire [2:0] L2BroadcastHub_1_io_outer_grant_bits_addr_beat;
  wire [2:0] L2BroadcastHub_1_io_outer_grant_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] L2BroadcastHub_1_io_outer_grant_bits_g_type;
  wire [63:0] L2BroadcastHub_1_io_outer_grant_bits_data;
  wire  L2BroadcastHub_1_io_outer_grant_bits_manager_id;
  wire  L2BroadcastHub_1_io_outer_finish_ready;
  wire  L2BroadcastHub_1_io_outer_finish_valid;
  wire  L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_outer_finish_bits_manager_id;
  wire  mmioManager_clk;
  wire  mmioManager_reset;
  wire  mmioManager_io_inner_acquire_ready;
  wire  mmioManager_io_inner_acquire_valid;
  wire [25:0] mmioManager_io_inner_acquire_bits_addr_block;
  wire [1:0] mmioManager_io_inner_acquire_bits_client_xact_id;
  wire [2:0] mmioManager_io_inner_acquire_bits_addr_beat;
  wire  mmioManager_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] mmioManager_io_inner_acquire_bits_a_type;
  wire [11:0] mmioManager_io_inner_acquire_bits_union;
  wire [63:0] mmioManager_io_inner_acquire_bits_data;
  wire  mmioManager_io_inner_acquire_bits_client_id;
  wire  mmioManager_io_inner_grant_ready;
  wire  mmioManager_io_inner_grant_valid;
  wire [2:0] mmioManager_io_inner_grant_bits_addr_beat;
  wire [1:0] mmioManager_io_inner_grant_bits_client_xact_id;
  wire [2:0] mmioManager_io_inner_grant_bits_manager_xact_id;
  wire  mmioManager_io_inner_grant_bits_is_builtin_type;
  wire [3:0] mmioManager_io_inner_grant_bits_g_type;
  wire [63:0] mmioManager_io_inner_grant_bits_data;
  wire  mmioManager_io_inner_grant_bits_client_id;
  wire  mmioManager_io_inner_finish_ready;
  wire  mmioManager_io_inner_finish_valid;
  wire [2:0] mmioManager_io_inner_finish_bits_manager_xact_id;
  wire  mmioManager_io_inner_probe_ready;
  wire  mmioManager_io_inner_probe_valid;
  wire [25:0] mmioManager_io_inner_probe_bits_addr_block;
  wire [1:0] mmioManager_io_inner_probe_bits_p_type;
  wire  mmioManager_io_inner_probe_bits_client_id;
  wire  mmioManager_io_inner_release_ready;
  wire  mmioManager_io_inner_release_valid;
  wire [2:0] mmioManager_io_inner_release_bits_addr_beat;
  wire [25:0] mmioManager_io_inner_release_bits_addr_block;
  wire [1:0] mmioManager_io_inner_release_bits_client_xact_id;
  wire  mmioManager_io_inner_release_bits_voluntary;
  wire [2:0] mmioManager_io_inner_release_bits_r_type;
  wire [63:0] mmioManager_io_inner_release_bits_data;
  wire  mmioManager_io_inner_release_bits_client_id;
  wire  mmioManager_io_incoherent_0;
  wire  mmioManager_io_outer_acquire_ready;
  wire  mmioManager_io_outer_acquire_valid;
  wire [25:0] mmioManager_io_outer_acquire_bits_addr_block;
  wire [1:0] mmioManager_io_outer_acquire_bits_client_xact_id;
  wire [2:0] mmioManager_io_outer_acquire_bits_addr_beat;
  wire  mmioManager_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] mmioManager_io_outer_acquire_bits_a_type;
  wire [11:0] mmioManager_io_outer_acquire_bits_union;
  wire [63:0] mmioManager_io_outer_acquire_bits_data;
  wire  mmioManager_io_outer_grant_ready;
  wire  mmioManager_io_outer_grant_valid;
  wire [2:0] mmioManager_io_outer_grant_bits_addr_beat;
  wire [1:0] mmioManager_io_outer_grant_bits_client_xact_id;
  wire  mmioManager_io_outer_grant_bits_manager_xact_id;
  wire  mmioManager_io_outer_grant_bits_is_builtin_type;
  wire [3:0] mmioManager_io_outer_grant_bits_g_type;
  wire [63:0] mmioManager_io_outer_grant_bits_data;
  wire  mem_ic_clk;
  wire  mem_ic_reset;
  wire  mem_ic_io_in_0_acquire_ready;
  wire  mem_ic_io_in_0_acquire_valid;
  wire [25:0] mem_ic_io_in_0_acquire_bits_addr_block;
  wire [2:0] mem_ic_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] mem_ic_io_in_0_acquire_bits_addr_beat;
  wire  mem_ic_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] mem_ic_io_in_0_acquire_bits_a_type;
  wire [11:0] mem_ic_io_in_0_acquire_bits_union;
  wire [63:0] mem_ic_io_in_0_acquire_bits_data;
  wire  mem_ic_io_in_0_grant_ready;
  wire  mem_ic_io_in_0_grant_valid;
  wire [2:0] mem_ic_io_in_0_grant_bits_addr_beat;
  wire [2:0] mem_ic_io_in_0_grant_bits_client_xact_id;
  wire  mem_ic_io_in_0_grant_bits_manager_xact_id;
  wire  mem_ic_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] mem_ic_io_in_0_grant_bits_g_type;
  wire [63:0] mem_ic_io_in_0_grant_bits_data;
  wire  mem_ic_io_out_0_acquire_ready;
  wire  mem_ic_io_out_0_acquire_valid;
  wire [25:0] mem_ic_io_out_0_acquire_bits_addr_block;
  wire [2:0] mem_ic_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] mem_ic_io_out_0_acquire_bits_addr_beat;
  wire  mem_ic_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] mem_ic_io_out_0_acquire_bits_a_type;
  wire [11:0] mem_ic_io_out_0_acquire_bits_union;
  wire [63:0] mem_ic_io_out_0_acquire_bits_data;
  wire  mem_ic_io_out_0_grant_ready;
  wire  mem_ic_io_out_0_grant_valid;
  wire [2:0] mem_ic_io_out_0_grant_bits_addr_beat;
  wire [2:0] mem_ic_io_out_0_grant_bits_client_xact_id;
  wire  mem_ic_io_out_0_grant_bits_manager_xact_id;
  wire  mem_ic_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] mem_ic_io_out_0_grant_bits_g_type;
  wire [63:0] mem_ic_io_out_0_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_clk;
  wire  ClientTileLinkIOUnwrapper_1_reset;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type;
  wire [11:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_probe_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_probe_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_valid;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type;
  wire [11:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_clk;
  wire  ClientTileLinkEnqueuer_1_reset;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type;
  wire [11:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_probe_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_valid;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  wire [11:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_probe_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_valid;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id;
  wire  NastiIOTileLinkIOConverter_1_clk;
  wire  NastiIOTileLinkIOConverter_1_reset;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_ready;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_valid;
  wire [25:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type;
  wire [11:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_ready;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_valid;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_valid;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user;
  wire  Queue_15_1_clk;
  wire  Queue_15_1_reset;
  wire  Queue_15_1_io_enq_ready;
  wire  Queue_15_1_io_enq_valid;
  wire [31:0] Queue_15_1_io_enq_bits_addr;
  wire [7:0] Queue_15_1_io_enq_bits_len;
  wire [2:0] Queue_15_1_io_enq_bits_size;
  wire [1:0] Queue_15_1_io_enq_bits_burst;
  wire  Queue_15_1_io_enq_bits_lock;
  wire [3:0] Queue_15_1_io_enq_bits_cache;
  wire [2:0] Queue_15_1_io_enq_bits_prot;
  wire [3:0] Queue_15_1_io_enq_bits_qos;
  wire [3:0] Queue_15_1_io_enq_bits_region;
  wire [4:0] Queue_15_1_io_enq_bits_id;
  wire  Queue_15_1_io_enq_bits_user;
  wire  Queue_15_1_io_deq_ready;
  wire  Queue_15_1_io_deq_valid;
  wire [31:0] Queue_15_1_io_deq_bits_addr;
  wire [7:0] Queue_15_1_io_deq_bits_len;
  wire [2:0] Queue_15_1_io_deq_bits_size;
  wire [1:0] Queue_15_1_io_deq_bits_burst;
  wire  Queue_15_1_io_deq_bits_lock;
  wire [3:0] Queue_15_1_io_deq_bits_cache;
  wire [2:0] Queue_15_1_io_deq_bits_prot;
  wire [3:0] Queue_15_1_io_deq_bits_qos;
  wire [3:0] Queue_15_1_io_deq_bits_region;
  wire [4:0] Queue_15_1_io_deq_bits_id;
  wire  Queue_15_1_io_deq_bits_user;
  wire  Queue_15_1_io_count;
  wire  Queue_16_1_clk;
  wire  Queue_16_1_reset;
  wire  Queue_16_1_io_enq_ready;
  wire  Queue_16_1_io_enq_valid;
  wire [31:0] Queue_16_1_io_enq_bits_addr;
  wire [7:0] Queue_16_1_io_enq_bits_len;
  wire [2:0] Queue_16_1_io_enq_bits_size;
  wire [1:0] Queue_16_1_io_enq_bits_burst;
  wire  Queue_16_1_io_enq_bits_lock;
  wire [3:0] Queue_16_1_io_enq_bits_cache;
  wire [2:0] Queue_16_1_io_enq_bits_prot;
  wire [3:0] Queue_16_1_io_enq_bits_qos;
  wire [3:0] Queue_16_1_io_enq_bits_region;
  wire [4:0] Queue_16_1_io_enq_bits_id;
  wire  Queue_16_1_io_enq_bits_user;
  wire  Queue_16_1_io_deq_ready;
  wire  Queue_16_1_io_deq_valid;
  wire [31:0] Queue_16_1_io_deq_bits_addr;
  wire [7:0] Queue_16_1_io_deq_bits_len;
  wire [2:0] Queue_16_1_io_deq_bits_size;
  wire [1:0] Queue_16_1_io_deq_bits_burst;
  wire  Queue_16_1_io_deq_bits_lock;
  wire [3:0] Queue_16_1_io_deq_bits_cache;
  wire [2:0] Queue_16_1_io_deq_bits_prot;
  wire [3:0] Queue_16_1_io_deq_bits_qos;
  wire [3:0] Queue_16_1_io_deq_bits_region;
  wire [4:0] Queue_16_1_io_deq_bits_id;
  wire  Queue_16_1_io_deq_bits_user;
  wire  Queue_16_1_io_count;
  wire  Queue_17_1_clk;
  wire  Queue_17_1_reset;
  wire  Queue_17_1_io_enq_ready;
  wire  Queue_17_1_io_enq_valid;
  wire [63:0] Queue_17_1_io_enq_bits_data;
  wire  Queue_17_1_io_enq_bits_last;
  wire [4:0] Queue_17_1_io_enq_bits_id;
  wire [7:0] Queue_17_1_io_enq_bits_strb;
  wire  Queue_17_1_io_enq_bits_user;
  wire  Queue_17_1_io_deq_ready;
  wire  Queue_17_1_io_deq_valid;
  wire [63:0] Queue_17_1_io_deq_bits_data;
  wire  Queue_17_1_io_deq_bits_last;
  wire [4:0] Queue_17_1_io_deq_bits_id;
  wire [7:0] Queue_17_1_io_deq_bits_strb;
  wire  Queue_17_1_io_deq_bits_user;
  wire [1:0] Queue_17_1_io_count;
  wire  Queue_18_1_clk;
  wire  Queue_18_1_reset;
  wire  Queue_18_1_io_enq_ready;
  wire  Queue_18_1_io_enq_valid;
  wire [1:0] Queue_18_1_io_enq_bits_resp;
  wire [63:0] Queue_18_1_io_enq_bits_data;
  wire  Queue_18_1_io_enq_bits_last;
  wire [4:0] Queue_18_1_io_enq_bits_id;
  wire  Queue_18_1_io_enq_bits_user;
  wire  Queue_18_1_io_deq_ready;
  wire  Queue_18_1_io_deq_valid;
  wire [1:0] Queue_18_1_io_deq_bits_resp;
  wire [63:0] Queue_18_1_io_deq_bits_data;
  wire  Queue_18_1_io_deq_bits_last;
  wire [4:0] Queue_18_1_io_deq_bits_id;
  wire  Queue_18_1_io_deq_bits_user;
  wire [1:0] Queue_18_1_io_count;
  wire  Queue_19_1_clk;
  wire  Queue_19_1_reset;
  wire  Queue_19_1_io_enq_ready;
  wire  Queue_19_1_io_enq_valid;
  wire [1:0] Queue_19_1_io_enq_bits_resp;
  wire [4:0] Queue_19_1_io_enq_bits_id;
  wire  Queue_19_1_io_enq_bits_user;
  wire  Queue_19_1_io_deq_ready;
  wire  Queue_19_1_io_deq_valid;
  wire [1:0] Queue_19_1_io_deq_bits_resp;
  wire [4:0] Queue_19_1_io_deq_bits_id;
  wire  Queue_19_1_io_deq_bits_user;
  wire  Queue_19_1_io_count;
  reg  GEN_0;
  reg [31:0] GEN_1;
  PortedTileLinkCrossbar l1tol2net (
    .clk(l1tol2net_clk),
    .reset(l1tol2net_reset),
    .io_clients_cached_0_acquire_ready(l1tol2net_io_clients_cached_0_acquire_ready),
    .io_clients_cached_0_acquire_valid(l1tol2net_io_clients_cached_0_acquire_valid),
    .io_clients_cached_0_acquire_bits_addr_block(l1tol2net_io_clients_cached_0_acquire_bits_addr_block),
    .io_clients_cached_0_acquire_bits_client_xact_id(l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id),
    .io_clients_cached_0_acquire_bits_addr_beat(l1tol2net_io_clients_cached_0_acquire_bits_addr_beat),
    .io_clients_cached_0_acquire_bits_is_builtin_type(l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type),
    .io_clients_cached_0_acquire_bits_a_type(l1tol2net_io_clients_cached_0_acquire_bits_a_type),
    .io_clients_cached_0_acquire_bits_union(l1tol2net_io_clients_cached_0_acquire_bits_union),
    .io_clients_cached_0_acquire_bits_data(l1tol2net_io_clients_cached_0_acquire_bits_data),
    .io_clients_cached_0_probe_ready(l1tol2net_io_clients_cached_0_probe_ready),
    .io_clients_cached_0_probe_valid(l1tol2net_io_clients_cached_0_probe_valid),
    .io_clients_cached_0_probe_bits_addr_block(l1tol2net_io_clients_cached_0_probe_bits_addr_block),
    .io_clients_cached_0_probe_bits_p_type(l1tol2net_io_clients_cached_0_probe_bits_p_type),
    .io_clients_cached_0_release_ready(l1tol2net_io_clients_cached_0_release_ready),
    .io_clients_cached_0_release_valid(l1tol2net_io_clients_cached_0_release_valid),
    .io_clients_cached_0_release_bits_addr_beat(l1tol2net_io_clients_cached_0_release_bits_addr_beat),
    .io_clients_cached_0_release_bits_addr_block(l1tol2net_io_clients_cached_0_release_bits_addr_block),
    .io_clients_cached_0_release_bits_client_xact_id(l1tol2net_io_clients_cached_0_release_bits_client_xact_id),
    .io_clients_cached_0_release_bits_voluntary(l1tol2net_io_clients_cached_0_release_bits_voluntary),
    .io_clients_cached_0_release_bits_r_type(l1tol2net_io_clients_cached_0_release_bits_r_type),
    .io_clients_cached_0_release_bits_data(l1tol2net_io_clients_cached_0_release_bits_data),
    .io_clients_cached_0_grant_ready(l1tol2net_io_clients_cached_0_grant_ready),
    .io_clients_cached_0_grant_valid(l1tol2net_io_clients_cached_0_grant_valid),
    .io_clients_cached_0_grant_bits_addr_beat(l1tol2net_io_clients_cached_0_grant_bits_addr_beat),
    .io_clients_cached_0_grant_bits_client_xact_id(l1tol2net_io_clients_cached_0_grant_bits_client_xact_id),
    .io_clients_cached_0_grant_bits_manager_xact_id(l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id),
    .io_clients_cached_0_grant_bits_is_builtin_type(l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type),
    .io_clients_cached_0_grant_bits_g_type(l1tol2net_io_clients_cached_0_grant_bits_g_type),
    .io_clients_cached_0_grant_bits_data(l1tol2net_io_clients_cached_0_grant_bits_data),
    .io_clients_cached_0_grant_bits_manager_id(l1tol2net_io_clients_cached_0_grant_bits_manager_id),
    .io_clients_cached_0_finish_ready(l1tol2net_io_clients_cached_0_finish_ready),
    .io_clients_cached_0_finish_valid(l1tol2net_io_clients_cached_0_finish_valid),
    .io_clients_cached_0_finish_bits_manager_xact_id(l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id),
    .io_clients_cached_0_finish_bits_manager_id(l1tol2net_io_clients_cached_0_finish_bits_manager_id),
    .io_clients_uncached_0_acquire_ready(l1tol2net_io_clients_uncached_0_acquire_ready),
    .io_clients_uncached_0_acquire_valid(l1tol2net_io_clients_uncached_0_acquire_valid),
    .io_clients_uncached_0_acquire_bits_addr_block(l1tol2net_io_clients_uncached_0_acquire_bits_addr_block),
    .io_clients_uncached_0_acquire_bits_client_xact_id(l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id),
    .io_clients_uncached_0_acquire_bits_addr_beat(l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat),
    .io_clients_uncached_0_acquire_bits_is_builtin_type(l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type),
    .io_clients_uncached_0_acquire_bits_a_type(l1tol2net_io_clients_uncached_0_acquire_bits_a_type),
    .io_clients_uncached_0_acquire_bits_union(l1tol2net_io_clients_uncached_0_acquire_bits_union),
    .io_clients_uncached_0_acquire_bits_data(l1tol2net_io_clients_uncached_0_acquire_bits_data),
    .io_clients_uncached_0_grant_ready(l1tol2net_io_clients_uncached_0_grant_ready),
    .io_clients_uncached_0_grant_valid(l1tol2net_io_clients_uncached_0_grant_valid),
    .io_clients_uncached_0_grant_bits_addr_beat(l1tol2net_io_clients_uncached_0_grant_bits_addr_beat),
    .io_clients_uncached_0_grant_bits_client_xact_id(l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id),
    .io_clients_uncached_0_grant_bits_manager_xact_id(l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id),
    .io_clients_uncached_0_grant_bits_is_builtin_type(l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type),
    .io_clients_uncached_0_grant_bits_g_type(l1tol2net_io_clients_uncached_0_grant_bits_g_type),
    .io_clients_uncached_0_grant_bits_data(l1tol2net_io_clients_uncached_0_grant_bits_data),
    .io_managers_0_acquire_ready(l1tol2net_io_managers_0_acquire_ready),
    .io_managers_0_acquire_valid(l1tol2net_io_managers_0_acquire_valid),
    .io_managers_0_acquire_bits_addr_block(l1tol2net_io_managers_0_acquire_bits_addr_block),
    .io_managers_0_acquire_bits_client_xact_id(l1tol2net_io_managers_0_acquire_bits_client_xact_id),
    .io_managers_0_acquire_bits_addr_beat(l1tol2net_io_managers_0_acquire_bits_addr_beat),
    .io_managers_0_acquire_bits_is_builtin_type(l1tol2net_io_managers_0_acquire_bits_is_builtin_type),
    .io_managers_0_acquire_bits_a_type(l1tol2net_io_managers_0_acquire_bits_a_type),
    .io_managers_0_acquire_bits_union(l1tol2net_io_managers_0_acquire_bits_union),
    .io_managers_0_acquire_bits_data(l1tol2net_io_managers_0_acquire_bits_data),
    .io_managers_0_acquire_bits_client_id(l1tol2net_io_managers_0_acquire_bits_client_id),
    .io_managers_0_grant_ready(l1tol2net_io_managers_0_grant_ready),
    .io_managers_0_grant_valid(l1tol2net_io_managers_0_grant_valid),
    .io_managers_0_grant_bits_addr_beat(l1tol2net_io_managers_0_grant_bits_addr_beat),
    .io_managers_0_grant_bits_client_xact_id(l1tol2net_io_managers_0_grant_bits_client_xact_id),
    .io_managers_0_grant_bits_manager_xact_id(l1tol2net_io_managers_0_grant_bits_manager_xact_id),
    .io_managers_0_grant_bits_is_builtin_type(l1tol2net_io_managers_0_grant_bits_is_builtin_type),
    .io_managers_0_grant_bits_g_type(l1tol2net_io_managers_0_grant_bits_g_type),
    .io_managers_0_grant_bits_data(l1tol2net_io_managers_0_grant_bits_data),
    .io_managers_0_grant_bits_client_id(l1tol2net_io_managers_0_grant_bits_client_id),
    .io_managers_0_finish_ready(l1tol2net_io_managers_0_finish_ready),
    .io_managers_0_finish_valid(l1tol2net_io_managers_0_finish_valid),
    .io_managers_0_finish_bits_manager_xact_id(l1tol2net_io_managers_0_finish_bits_manager_xact_id),
    .io_managers_0_probe_ready(l1tol2net_io_managers_0_probe_ready),
    .io_managers_0_probe_valid(l1tol2net_io_managers_0_probe_valid),
    .io_managers_0_probe_bits_addr_block(l1tol2net_io_managers_0_probe_bits_addr_block),
    .io_managers_0_probe_bits_p_type(l1tol2net_io_managers_0_probe_bits_p_type),
    .io_managers_0_probe_bits_client_id(l1tol2net_io_managers_0_probe_bits_client_id),
    .io_managers_0_release_ready(l1tol2net_io_managers_0_release_ready),
    .io_managers_0_release_valid(l1tol2net_io_managers_0_release_valid),
    .io_managers_0_release_bits_addr_beat(l1tol2net_io_managers_0_release_bits_addr_beat),
    .io_managers_0_release_bits_addr_block(l1tol2net_io_managers_0_release_bits_addr_block),
    .io_managers_0_release_bits_client_xact_id(l1tol2net_io_managers_0_release_bits_client_xact_id),
    .io_managers_0_release_bits_voluntary(l1tol2net_io_managers_0_release_bits_voluntary),
    .io_managers_0_release_bits_r_type(l1tol2net_io_managers_0_release_bits_r_type),
    .io_managers_0_release_bits_data(l1tol2net_io_managers_0_release_bits_data),
    .io_managers_0_release_bits_client_id(l1tol2net_io_managers_0_release_bits_client_id),
    .io_managers_1_acquire_ready(l1tol2net_io_managers_1_acquire_ready),
    .io_managers_1_acquire_valid(l1tol2net_io_managers_1_acquire_valid),
    .io_managers_1_acquire_bits_addr_block(l1tol2net_io_managers_1_acquire_bits_addr_block),
    .io_managers_1_acquire_bits_client_xact_id(l1tol2net_io_managers_1_acquire_bits_client_xact_id),
    .io_managers_1_acquire_bits_addr_beat(l1tol2net_io_managers_1_acquire_bits_addr_beat),
    .io_managers_1_acquire_bits_is_builtin_type(l1tol2net_io_managers_1_acquire_bits_is_builtin_type),
    .io_managers_1_acquire_bits_a_type(l1tol2net_io_managers_1_acquire_bits_a_type),
    .io_managers_1_acquire_bits_union(l1tol2net_io_managers_1_acquire_bits_union),
    .io_managers_1_acquire_bits_data(l1tol2net_io_managers_1_acquire_bits_data),
    .io_managers_1_acquire_bits_client_id(l1tol2net_io_managers_1_acquire_bits_client_id),
    .io_managers_1_grant_ready(l1tol2net_io_managers_1_grant_ready),
    .io_managers_1_grant_valid(l1tol2net_io_managers_1_grant_valid),
    .io_managers_1_grant_bits_addr_beat(l1tol2net_io_managers_1_grant_bits_addr_beat),
    .io_managers_1_grant_bits_client_xact_id(l1tol2net_io_managers_1_grant_bits_client_xact_id),
    .io_managers_1_grant_bits_manager_xact_id(l1tol2net_io_managers_1_grant_bits_manager_xact_id),
    .io_managers_1_grant_bits_is_builtin_type(l1tol2net_io_managers_1_grant_bits_is_builtin_type),
    .io_managers_1_grant_bits_g_type(l1tol2net_io_managers_1_grant_bits_g_type),
    .io_managers_1_grant_bits_data(l1tol2net_io_managers_1_grant_bits_data),
    .io_managers_1_grant_bits_client_id(l1tol2net_io_managers_1_grant_bits_client_id),
    .io_managers_1_finish_ready(l1tol2net_io_managers_1_finish_ready),
    .io_managers_1_finish_valid(l1tol2net_io_managers_1_finish_valid),
    .io_managers_1_finish_bits_manager_xact_id(l1tol2net_io_managers_1_finish_bits_manager_xact_id),
    .io_managers_1_probe_ready(l1tol2net_io_managers_1_probe_ready),
    .io_managers_1_probe_valid(l1tol2net_io_managers_1_probe_valid),
    .io_managers_1_probe_bits_addr_block(l1tol2net_io_managers_1_probe_bits_addr_block),
    .io_managers_1_probe_bits_p_type(l1tol2net_io_managers_1_probe_bits_p_type),
    .io_managers_1_probe_bits_client_id(l1tol2net_io_managers_1_probe_bits_client_id),
    .io_managers_1_release_ready(l1tol2net_io_managers_1_release_ready),
    .io_managers_1_release_valid(l1tol2net_io_managers_1_release_valid),
    .io_managers_1_release_bits_addr_beat(l1tol2net_io_managers_1_release_bits_addr_beat),
    .io_managers_1_release_bits_addr_block(l1tol2net_io_managers_1_release_bits_addr_block),
    .io_managers_1_release_bits_client_xact_id(l1tol2net_io_managers_1_release_bits_client_xact_id),
    .io_managers_1_release_bits_voluntary(l1tol2net_io_managers_1_release_bits_voluntary),
    .io_managers_1_release_bits_r_type(l1tol2net_io_managers_1_release_bits_r_type),
    .io_managers_1_release_bits_data(l1tol2net_io_managers_1_release_bits_data),
    .io_managers_1_release_bits_client_id(l1tol2net_io_managers_1_release_bits_client_id)
  );
  L2BroadcastHub L2BroadcastHub_1 (
    .clk(L2BroadcastHub_1_clk),
    .reset(L2BroadcastHub_1_reset),
    .io_inner_acquire_ready(L2BroadcastHub_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(L2BroadcastHub_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(L2BroadcastHub_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(L2BroadcastHub_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(L2BroadcastHub_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(L2BroadcastHub_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(L2BroadcastHub_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(L2BroadcastHub_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(L2BroadcastHub_1_io_inner_grant_ready),
    .io_inner_grant_valid(L2BroadcastHub_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(L2BroadcastHub_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(L2BroadcastHub_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(L2BroadcastHub_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(L2BroadcastHub_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(L2BroadcastHub_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(L2BroadcastHub_1_io_inner_finish_ready),
    .io_inner_finish_valid(L2BroadcastHub_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(L2BroadcastHub_1_io_inner_probe_ready),
    .io_inner_probe_valid(L2BroadcastHub_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(L2BroadcastHub_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(L2BroadcastHub_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(L2BroadcastHub_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(L2BroadcastHub_1_io_inner_release_ready),
    .io_inner_release_valid(L2BroadcastHub_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(L2BroadcastHub_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(L2BroadcastHub_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(L2BroadcastHub_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(L2BroadcastHub_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(L2BroadcastHub_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(L2BroadcastHub_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(L2BroadcastHub_1_io_inner_release_bits_client_id),
    .io_incoherent_0(L2BroadcastHub_1_io_incoherent_0),
    .io_outer_acquire_ready(L2BroadcastHub_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(L2BroadcastHub_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(L2BroadcastHub_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(L2BroadcastHub_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(L2BroadcastHub_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(L2BroadcastHub_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(L2BroadcastHub_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(L2BroadcastHub_1_io_outer_probe_ready),
    .io_outer_probe_valid(L2BroadcastHub_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(L2BroadcastHub_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(L2BroadcastHub_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(L2BroadcastHub_1_io_outer_release_ready),
    .io_outer_release_valid(L2BroadcastHub_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(L2BroadcastHub_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(L2BroadcastHub_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(L2BroadcastHub_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(L2BroadcastHub_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(L2BroadcastHub_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(L2BroadcastHub_1_io_outer_release_bits_data),
    .io_outer_grant_ready(L2BroadcastHub_1_io_outer_grant_ready),
    .io_outer_grant_valid(L2BroadcastHub_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(L2BroadcastHub_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(L2BroadcastHub_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(L2BroadcastHub_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(L2BroadcastHub_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(L2BroadcastHub_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(L2BroadcastHub_1_io_outer_finish_ready),
    .io_outer_finish_valid(L2BroadcastHub_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(L2BroadcastHub_1_io_outer_finish_bits_manager_id)
  );
  MMIOTileLinkManager mmioManager (
    .clk(mmioManager_clk),
    .reset(mmioManager_reset),
    .io_inner_acquire_ready(mmioManager_io_inner_acquire_ready),
    .io_inner_acquire_valid(mmioManager_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(mmioManager_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(mmioManager_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(mmioManager_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(mmioManager_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(mmioManager_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(mmioManager_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(mmioManager_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(mmioManager_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(mmioManager_io_inner_grant_ready),
    .io_inner_grant_valid(mmioManager_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(mmioManager_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(mmioManager_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(mmioManager_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(mmioManager_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(mmioManager_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(mmioManager_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(mmioManager_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(mmioManager_io_inner_finish_ready),
    .io_inner_finish_valid(mmioManager_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(mmioManager_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(mmioManager_io_inner_probe_ready),
    .io_inner_probe_valid(mmioManager_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(mmioManager_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(mmioManager_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(mmioManager_io_inner_probe_bits_client_id),
    .io_inner_release_ready(mmioManager_io_inner_release_ready),
    .io_inner_release_valid(mmioManager_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(mmioManager_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(mmioManager_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(mmioManager_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(mmioManager_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(mmioManager_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(mmioManager_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(mmioManager_io_inner_release_bits_client_id),
    .io_incoherent_0(mmioManager_io_incoherent_0),
    .io_outer_acquire_ready(mmioManager_io_outer_acquire_ready),
    .io_outer_acquire_valid(mmioManager_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(mmioManager_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(mmioManager_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(mmioManager_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(mmioManager_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(mmioManager_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(mmioManager_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(mmioManager_io_outer_acquire_bits_data),
    .io_outer_grant_ready(mmioManager_io_outer_grant_ready),
    .io_outer_grant_valid(mmioManager_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(mmioManager_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(mmioManager_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(mmioManager_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(mmioManager_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(mmioManager_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(mmioManager_io_outer_grant_bits_data)
  );
  TileLinkMemoryInterconnect mem_ic (
    .clk(mem_ic_clk),
    .reset(mem_ic_reset),
    .io_in_0_acquire_ready(mem_ic_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(mem_ic_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(mem_ic_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(mem_ic_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(mem_ic_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(mem_ic_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(mem_ic_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(mem_ic_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(mem_ic_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(mem_ic_io_in_0_grant_ready),
    .io_in_0_grant_valid(mem_ic_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(mem_ic_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(mem_ic_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(mem_ic_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(mem_ic_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(mem_ic_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(mem_ic_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(mem_ic_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(mem_ic_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(mem_ic_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(mem_ic_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(mem_ic_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(mem_ic_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(mem_ic_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(mem_ic_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(mem_ic_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(mem_ic_io_out_0_grant_ready),
    .io_out_0_grant_valid(mem_ic_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(mem_ic_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(mem_ic_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(mem_ic_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(mem_ic_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(mem_ic_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(mem_ic_io_out_0_grant_bits_data)
  );
  ClientTileLinkIOUnwrapper ClientTileLinkIOUnwrapper_1 (
    .clk(ClientTileLinkIOUnwrapper_1_clk),
    .reset(ClientTileLinkIOUnwrapper_1_reset),
    .io_in_acquire_ready(ClientTileLinkIOUnwrapper_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientTileLinkIOUnwrapper_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data),
    .io_in_probe_ready(ClientTileLinkIOUnwrapper_1_io_in_probe_ready),
    .io_in_probe_valid(ClientTileLinkIOUnwrapper_1_io_in_probe_valid),
    .io_in_probe_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block),
    .io_in_probe_bits_p_type(ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type),
    .io_in_release_ready(ClientTileLinkIOUnwrapper_1_io_in_release_ready),
    .io_in_release_valid(ClientTileLinkIOUnwrapper_1_io_in_release_valid),
    .io_in_release_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat),
    .io_in_release_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block),
    .io_in_release_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id),
    .io_in_release_bits_voluntary(ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary),
    .io_in_release_bits_r_type(ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type),
    .io_in_release_bits_data(ClientTileLinkIOUnwrapper_1_io_in_release_bits_data),
    .io_in_grant_ready(ClientTileLinkIOUnwrapper_1_io_in_grant_ready),
    .io_in_grant_valid(ClientTileLinkIOUnwrapper_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data),
    .io_in_grant_bits_manager_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id),
    .io_in_finish_ready(ClientTileLinkIOUnwrapper_1_io_in_finish_ready),
    .io_in_finish_valid(ClientTileLinkIOUnwrapper_1_io_in_finish_valid),
    .io_in_finish_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id),
    .io_in_finish_bits_manager_id(ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id),
    .io_out_acquire_ready(ClientTileLinkIOUnwrapper_1_io_out_acquire_ready),
    .io_out_acquire_valid(ClientTileLinkIOUnwrapper_1_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientTileLinkIOUnwrapper_1_io_out_grant_ready),
    .io_out_grant_valid(ClientTileLinkIOUnwrapper_1_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data)
  );
  ClientTileLinkEnqueuer ClientTileLinkEnqueuer_1 (
    .clk(ClientTileLinkEnqueuer_1_clk),
    .reset(ClientTileLinkEnqueuer_1_reset),
    .io_inner_acquire_ready(ClientTileLinkEnqueuer_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(ClientTileLinkEnqueuer_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data),
    .io_inner_probe_ready(ClientTileLinkEnqueuer_1_io_inner_probe_ready),
    .io_inner_probe_valid(ClientTileLinkEnqueuer_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type),
    .io_inner_release_ready(ClientTileLinkEnqueuer_1_io_inner_release_ready),
    .io_inner_release_valid(ClientTileLinkEnqueuer_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(ClientTileLinkEnqueuer_1_io_inner_release_bits_data),
    .io_inner_grant_ready(ClientTileLinkEnqueuer_1_io_inner_grant_ready),
    .io_inner_grant_valid(ClientTileLinkEnqueuer_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(ClientTileLinkEnqueuer_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_manager_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id),
    .io_inner_finish_ready(ClientTileLinkEnqueuer_1_io_inner_finish_ready),
    .io_inner_finish_valid(ClientTileLinkEnqueuer_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_finish_bits_manager_id(ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id),
    .io_outer_acquire_ready(ClientTileLinkEnqueuer_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(ClientTileLinkEnqueuer_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(ClientTileLinkEnqueuer_1_io_outer_probe_ready),
    .io_outer_probe_valid(ClientTileLinkEnqueuer_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(ClientTileLinkEnqueuer_1_io_outer_release_ready),
    .io_outer_release_valid(ClientTileLinkEnqueuer_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(ClientTileLinkEnqueuer_1_io_outer_release_bits_data),
    .io_outer_grant_ready(ClientTileLinkEnqueuer_1_io_outer_grant_ready),
    .io_outer_grant_valid(ClientTileLinkEnqueuer_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(ClientTileLinkEnqueuer_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(ClientTileLinkEnqueuer_1_io_outer_finish_ready),
    .io_outer_finish_valid(ClientTileLinkEnqueuer_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id)
  );
  NastiIOTileLinkIOConverter NastiIOTileLinkIOConverter_1 (
    .clk(NastiIOTileLinkIOConverter_1_clk),
    .reset(NastiIOTileLinkIOConverter_1_reset),
    .io_tl_acquire_ready(NastiIOTileLinkIOConverter_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(NastiIOTileLinkIOConverter_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(NastiIOTileLinkIOConverter_1_io_tl_grant_ready),
    .io_tl_grant_valid(NastiIOTileLinkIOConverter_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data),
    .io_nasti_aw_ready(NastiIOTileLinkIOConverter_1_io_nasti_aw_ready),
    .io_nasti_aw_valid(NastiIOTileLinkIOConverter_1_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user),
    .io_nasti_w_ready(NastiIOTileLinkIOConverter_1_io_nasti_w_ready),
    .io_nasti_w_valid(NastiIOTileLinkIOConverter_1_io_nasti_w_valid),
    .io_nasti_w_bits_data(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user),
    .io_nasti_b_ready(NastiIOTileLinkIOConverter_1_io_nasti_b_ready),
    .io_nasti_b_valid(NastiIOTileLinkIOConverter_1_io_nasti_b_valid),
    .io_nasti_b_bits_resp(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user),
    .io_nasti_ar_ready(NastiIOTileLinkIOConverter_1_io_nasti_ar_ready),
    .io_nasti_ar_valid(NastiIOTileLinkIOConverter_1_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user),
    .io_nasti_r_ready(NastiIOTileLinkIOConverter_1_io_nasti_r_ready),
    .io_nasti_r_valid(NastiIOTileLinkIOConverter_1_io_nasti_r_valid),
    .io_nasti_r_bits_resp(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user)
  );
  Queue_15 Queue_15_1 (
    .clk(Queue_15_1_clk),
    .reset(Queue_15_1_reset),
    .io_enq_ready(Queue_15_1_io_enq_ready),
    .io_enq_valid(Queue_15_1_io_enq_valid),
    .io_enq_bits_addr(Queue_15_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_15_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_15_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_15_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_15_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_15_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_15_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_15_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_15_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_15_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_15_1_io_enq_bits_user),
    .io_deq_ready(Queue_15_1_io_deq_ready),
    .io_deq_valid(Queue_15_1_io_deq_valid),
    .io_deq_bits_addr(Queue_15_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_15_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_15_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_15_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_15_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_15_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_15_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_15_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_15_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_15_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_15_1_io_deq_bits_user),
    .io_count(Queue_15_1_io_count)
  );
  Queue_15 Queue_16_1 (
    .clk(Queue_16_1_clk),
    .reset(Queue_16_1_reset),
    .io_enq_ready(Queue_16_1_io_enq_ready),
    .io_enq_valid(Queue_16_1_io_enq_valid),
    .io_enq_bits_addr(Queue_16_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_16_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_16_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_16_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_16_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_16_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_16_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_16_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_16_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_16_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_16_1_io_enq_bits_user),
    .io_deq_ready(Queue_16_1_io_deq_ready),
    .io_deq_valid(Queue_16_1_io_deq_valid),
    .io_deq_bits_addr(Queue_16_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_16_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_16_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_16_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_16_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_16_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_16_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_16_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_16_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_16_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_16_1_io_deq_bits_user),
    .io_count(Queue_16_1_io_count)
  );
  Queue_17 Queue_17_1 (
    .clk(Queue_17_1_clk),
    .reset(Queue_17_1_reset),
    .io_enq_ready(Queue_17_1_io_enq_ready),
    .io_enq_valid(Queue_17_1_io_enq_valid),
    .io_enq_bits_data(Queue_17_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_17_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_17_1_io_enq_bits_id),
    .io_enq_bits_strb(Queue_17_1_io_enq_bits_strb),
    .io_enq_bits_user(Queue_17_1_io_enq_bits_user),
    .io_deq_ready(Queue_17_1_io_deq_ready),
    .io_deq_valid(Queue_17_1_io_deq_valid),
    .io_deq_bits_data(Queue_17_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_17_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_17_1_io_deq_bits_id),
    .io_deq_bits_strb(Queue_17_1_io_deq_bits_strb),
    .io_deq_bits_user(Queue_17_1_io_deq_bits_user),
    .io_count(Queue_17_1_io_count)
  );
  Queue_18 Queue_18_1 (
    .clk(Queue_18_1_clk),
    .reset(Queue_18_1_reset),
    .io_enq_ready(Queue_18_1_io_enq_ready),
    .io_enq_valid(Queue_18_1_io_enq_valid),
    .io_enq_bits_resp(Queue_18_1_io_enq_bits_resp),
    .io_enq_bits_data(Queue_18_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_18_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_18_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_18_1_io_enq_bits_user),
    .io_deq_ready(Queue_18_1_io_deq_ready),
    .io_deq_valid(Queue_18_1_io_deq_valid),
    .io_deq_bits_resp(Queue_18_1_io_deq_bits_resp),
    .io_deq_bits_data(Queue_18_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_18_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_18_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_18_1_io_deq_bits_user),
    .io_count(Queue_18_1_io_count)
  );
  Queue_19 Queue_19_1 (
    .clk(Queue_19_1_clk),
    .reset(Queue_19_1_reset),
    .io_enq_ready(Queue_19_1_io_enq_ready),
    .io_enq_valid(Queue_19_1_io_enq_valid),
    .io_enq_bits_resp(Queue_19_1_io_enq_bits_resp),
    .io_enq_bits_id(Queue_19_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_19_1_io_enq_bits_user),
    .io_deq_ready(Queue_19_1_io_deq_ready),
    .io_deq_valid(Queue_19_1_io_deq_valid),
    .io_deq_bits_resp(Queue_19_1_io_deq_bits_resp),
    .io_deq_bits_id(Queue_19_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_19_1_io_deq_bits_user),
    .io_count(Queue_19_1_io_count)
  );
  assign io_tiles_cached_0_acquire_ready = l1tol2net_io_clients_cached_0_acquire_ready;
  assign io_tiles_cached_0_probe_valid = l1tol2net_io_clients_cached_0_probe_valid;
  assign io_tiles_cached_0_probe_bits_addr_block = l1tol2net_io_clients_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_bits_p_type = l1tol2net_io_clients_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_release_ready = l1tol2net_io_clients_cached_0_release_ready;
  assign io_tiles_cached_0_grant_valid = l1tol2net_io_clients_cached_0_grant_valid;
  assign io_tiles_cached_0_grant_bits_addr_beat = l1tol2net_io_clients_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_bits_client_xact_id = l1tol2net_io_clients_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_g_type = l1tol2net_io_clients_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_data = l1tol2net_io_clients_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_manager_id = l1tol2net_io_clients_cached_0_grant_bits_manager_id;
  assign io_tiles_cached_0_finish_ready = l1tol2net_io_clients_cached_0_finish_ready;
  assign io_tiles_uncached_0_acquire_ready = l1tol2net_io_clients_uncached_0_acquire_ready;
  assign io_tiles_uncached_0_grant_valid = l1tol2net_io_clients_uncached_0_grant_valid;
  assign io_tiles_uncached_0_grant_bits_addr_beat = l1tol2net_io_clients_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_g_type = l1tol2net_io_clients_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_data = l1tol2net_io_clients_uncached_0_grant_bits_data;
  assign io_mem_axi_0_aw_valid = Queue_16_1_io_deq_valid;
  assign io_mem_axi_0_aw_bits_addr = Queue_16_1_io_deq_bits_addr;
  assign io_mem_axi_0_aw_bits_len = Queue_16_1_io_deq_bits_len;
  assign io_mem_axi_0_aw_bits_size = Queue_16_1_io_deq_bits_size;
  assign io_mem_axi_0_aw_bits_burst = Queue_16_1_io_deq_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = Queue_16_1_io_deq_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = 4'h3;
  assign io_mem_axi_0_aw_bits_prot = Queue_16_1_io_deq_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = Queue_16_1_io_deq_bits_qos;
  assign io_mem_axi_0_aw_bits_region = Queue_16_1_io_deq_bits_region;
  assign io_mem_axi_0_aw_bits_id = Queue_16_1_io_deq_bits_id;
  assign io_mem_axi_0_aw_bits_user = Queue_16_1_io_deq_bits_user;
  assign io_mem_axi_0_w_valid = Queue_17_1_io_deq_valid;
  assign io_mem_axi_0_w_bits_data = Queue_17_1_io_deq_bits_data;
  assign io_mem_axi_0_w_bits_last = Queue_17_1_io_deq_bits_last;
  assign io_mem_axi_0_w_bits_id = Queue_17_1_io_deq_bits_id;
  assign io_mem_axi_0_w_bits_strb = Queue_17_1_io_deq_bits_strb;
  assign io_mem_axi_0_w_bits_user = Queue_17_1_io_deq_bits_user;
  assign io_mem_axi_0_b_ready = Queue_19_1_io_enq_ready;
  assign io_mem_axi_0_ar_valid = Queue_15_1_io_deq_valid;
  assign io_mem_axi_0_ar_bits_addr = Queue_15_1_io_deq_bits_addr;
  assign io_mem_axi_0_ar_bits_len = Queue_15_1_io_deq_bits_len;
  assign io_mem_axi_0_ar_bits_size = Queue_15_1_io_deq_bits_size;
  assign io_mem_axi_0_ar_bits_burst = Queue_15_1_io_deq_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = Queue_15_1_io_deq_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = 4'h3;
  assign io_mem_axi_0_ar_bits_prot = Queue_15_1_io_deq_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = Queue_15_1_io_deq_bits_qos;
  assign io_mem_axi_0_ar_bits_region = Queue_15_1_io_deq_bits_region;
  assign io_mem_axi_0_ar_bits_id = Queue_15_1_io_deq_bits_id;
  assign io_mem_axi_0_ar_bits_user = Queue_15_1_io_deq_bits_user;
  assign io_mem_axi_0_r_ready = Queue_18_1_io_enq_ready;
  assign io_mmio_acquire_valid = mmioManager_io_outer_acquire_valid;
  assign io_mmio_acquire_bits_addr_block = mmioManager_io_outer_acquire_bits_addr_block;
  assign io_mmio_acquire_bits_client_xact_id = mmioManager_io_outer_acquire_bits_client_xact_id;
  assign io_mmio_acquire_bits_addr_beat = mmioManager_io_outer_acquire_bits_addr_beat;
  assign io_mmio_acquire_bits_is_builtin_type = mmioManager_io_outer_acquire_bits_is_builtin_type;
  assign io_mmio_acquire_bits_a_type = mmioManager_io_outer_acquire_bits_a_type;
  assign io_mmio_acquire_bits_union = mmioManager_io_outer_acquire_bits_union;
  assign io_mmio_acquire_bits_data = mmioManager_io_outer_acquire_bits_data;
  assign io_mmio_grant_ready = mmioManager_io_outer_grant_ready;
  assign l1tol2net_clk = clk;
  assign l1tol2net_reset = reset;
  assign l1tol2net_io_clients_cached_0_acquire_valid = io_tiles_cached_0_acquire_valid;
  assign l1tol2net_io_clients_cached_0_acquire_bits_addr_block = io_tiles_cached_0_acquire_bits_addr_block;
  assign l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id = io_tiles_cached_0_acquire_bits_client_xact_id;
  assign l1tol2net_io_clients_cached_0_acquire_bits_addr_beat = io_tiles_cached_0_acquire_bits_addr_beat;
  assign l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type = io_tiles_cached_0_acquire_bits_is_builtin_type;
  assign l1tol2net_io_clients_cached_0_acquire_bits_a_type = io_tiles_cached_0_acquire_bits_a_type;
  assign l1tol2net_io_clients_cached_0_acquire_bits_union = io_tiles_cached_0_acquire_bits_union;
  assign l1tol2net_io_clients_cached_0_acquire_bits_data = io_tiles_cached_0_acquire_bits_data;
  assign l1tol2net_io_clients_cached_0_probe_ready = io_tiles_cached_0_probe_ready;
  assign l1tol2net_io_clients_cached_0_release_valid = io_tiles_cached_0_release_valid;
  assign l1tol2net_io_clients_cached_0_release_bits_addr_beat = io_tiles_cached_0_release_bits_addr_beat;
  assign l1tol2net_io_clients_cached_0_release_bits_addr_block = io_tiles_cached_0_release_bits_addr_block;
  assign l1tol2net_io_clients_cached_0_release_bits_client_xact_id = io_tiles_cached_0_release_bits_client_xact_id;
  assign l1tol2net_io_clients_cached_0_release_bits_voluntary = io_tiles_cached_0_release_bits_voluntary;
  assign l1tol2net_io_clients_cached_0_release_bits_r_type = io_tiles_cached_0_release_bits_r_type;
  assign l1tol2net_io_clients_cached_0_release_bits_data = io_tiles_cached_0_release_bits_data;
  assign l1tol2net_io_clients_cached_0_grant_ready = io_tiles_cached_0_grant_ready;
  assign l1tol2net_io_clients_cached_0_finish_valid = io_tiles_cached_0_finish_valid;
  assign l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id = io_tiles_cached_0_finish_bits_manager_xact_id;
  assign l1tol2net_io_clients_cached_0_finish_bits_manager_id = io_tiles_cached_0_finish_bits_manager_id;
  assign l1tol2net_io_clients_uncached_0_acquire_valid = io_tiles_uncached_0_acquire_valid;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_addr_block = io_tiles_uncached_0_acquire_bits_addr_block;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id = io_tiles_uncached_0_acquire_bits_client_xact_id;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat = io_tiles_uncached_0_acquire_bits_addr_beat;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type = io_tiles_uncached_0_acquire_bits_is_builtin_type;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_a_type = io_tiles_uncached_0_acquire_bits_a_type;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_union = io_tiles_uncached_0_acquire_bits_union;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_data = io_tiles_uncached_0_acquire_bits_data;
  assign l1tol2net_io_clients_uncached_0_grant_ready = io_tiles_uncached_0_grant_ready;
  assign l1tol2net_io_managers_0_acquire_ready = L2BroadcastHub_1_io_inner_acquire_ready;
  assign l1tol2net_io_managers_0_grant_valid = L2BroadcastHub_1_io_inner_grant_valid;
  assign l1tol2net_io_managers_0_grant_bits_addr_beat = L2BroadcastHub_1_io_inner_grant_bits_addr_beat;
  assign l1tol2net_io_managers_0_grant_bits_client_xact_id = L2BroadcastHub_1_io_inner_grant_bits_client_xact_id;
  assign l1tol2net_io_managers_0_grant_bits_manager_xact_id = L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id;
  assign l1tol2net_io_managers_0_grant_bits_is_builtin_type = L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type;
  assign l1tol2net_io_managers_0_grant_bits_g_type = L2BroadcastHub_1_io_inner_grant_bits_g_type;
  assign l1tol2net_io_managers_0_grant_bits_data = L2BroadcastHub_1_io_inner_grant_bits_data;
  assign l1tol2net_io_managers_0_grant_bits_client_id = L2BroadcastHub_1_io_inner_grant_bits_client_id;
  assign l1tol2net_io_managers_0_finish_ready = L2BroadcastHub_1_io_inner_finish_ready;
  assign l1tol2net_io_managers_0_probe_valid = L2BroadcastHub_1_io_inner_probe_valid;
  assign l1tol2net_io_managers_0_probe_bits_addr_block = L2BroadcastHub_1_io_inner_probe_bits_addr_block;
  assign l1tol2net_io_managers_0_probe_bits_p_type = L2BroadcastHub_1_io_inner_probe_bits_p_type;
  assign l1tol2net_io_managers_0_probe_bits_client_id = L2BroadcastHub_1_io_inner_probe_bits_client_id;
  assign l1tol2net_io_managers_0_release_ready = L2BroadcastHub_1_io_inner_release_ready;
  assign l1tol2net_io_managers_1_acquire_ready = mmioManager_io_inner_acquire_ready;
  assign l1tol2net_io_managers_1_grant_valid = mmioManager_io_inner_grant_valid;
  assign l1tol2net_io_managers_1_grant_bits_addr_beat = mmioManager_io_inner_grant_bits_addr_beat;
  assign l1tol2net_io_managers_1_grant_bits_client_xact_id = mmioManager_io_inner_grant_bits_client_xact_id;
  assign l1tol2net_io_managers_1_grant_bits_manager_xact_id = mmioManager_io_inner_grant_bits_manager_xact_id;
  assign l1tol2net_io_managers_1_grant_bits_is_builtin_type = mmioManager_io_inner_grant_bits_is_builtin_type;
  assign l1tol2net_io_managers_1_grant_bits_g_type = mmioManager_io_inner_grant_bits_g_type;
  assign l1tol2net_io_managers_1_grant_bits_data = mmioManager_io_inner_grant_bits_data;
  assign l1tol2net_io_managers_1_grant_bits_client_id = mmioManager_io_inner_grant_bits_client_id;
  assign l1tol2net_io_managers_1_finish_ready = mmioManager_io_inner_finish_ready;
  assign l1tol2net_io_managers_1_probe_valid = mmioManager_io_inner_probe_valid;
  assign l1tol2net_io_managers_1_probe_bits_addr_block = mmioManager_io_inner_probe_bits_addr_block;
  assign l1tol2net_io_managers_1_probe_bits_p_type = mmioManager_io_inner_probe_bits_p_type;
  assign l1tol2net_io_managers_1_probe_bits_client_id = mmioManager_io_inner_probe_bits_client_id;
  assign l1tol2net_io_managers_1_release_ready = mmioManager_io_inner_release_ready;
  assign L2BroadcastHub_1_clk = clk;
  assign L2BroadcastHub_1_reset = reset;
  assign L2BroadcastHub_1_io_inner_acquire_valid = l1tol2net_io_managers_0_acquire_valid;
  assign L2BroadcastHub_1_io_inner_acquire_bits_addr_block = l1tol2net_io_managers_0_acquire_bits_addr_block;
  assign L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id = l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  assign L2BroadcastHub_1_io_inner_acquire_bits_addr_beat = l1tol2net_io_managers_0_acquire_bits_addr_beat;
  assign L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type = l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  assign L2BroadcastHub_1_io_inner_acquire_bits_a_type = l1tol2net_io_managers_0_acquire_bits_a_type;
  assign L2BroadcastHub_1_io_inner_acquire_bits_union = l1tol2net_io_managers_0_acquire_bits_union;
  assign L2BroadcastHub_1_io_inner_acquire_bits_data = l1tol2net_io_managers_0_acquire_bits_data;
  assign L2BroadcastHub_1_io_inner_acquire_bits_client_id = l1tol2net_io_managers_0_acquire_bits_client_id;
  assign L2BroadcastHub_1_io_inner_grant_ready = l1tol2net_io_managers_0_grant_ready;
  assign L2BroadcastHub_1_io_inner_finish_valid = l1tol2net_io_managers_0_finish_valid;
  assign L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id = l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  assign L2BroadcastHub_1_io_inner_probe_ready = l1tol2net_io_managers_0_probe_ready;
  assign L2BroadcastHub_1_io_inner_release_valid = l1tol2net_io_managers_0_release_valid;
  assign L2BroadcastHub_1_io_inner_release_bits_addr_beat = l1tol2net_io_managers_0_release_bits_addr_beat;
  assign L2BroadcastHub_1_io_inner_release_bits_addr_block = l1tol2net_io_managers_0_release_bits_addr_block;
  assign L2BroadcastHub_1_io_inner_release_bits_client_xact_id = l1tol2net_io_managers_0_release_bits_client_xact_id;
  assign L2BroadcastHub_1_io_inner_release_bits_voluntary = l1tol2net_io_managers_0_release_bits_voluntary;
  assign L2BroadcastHub_1_io_inner_release_bits_r_type = l1tol2net_io_managers_0_release_bits_r_type;
  assign L2BroadcastHub_1_io_inner_release_bits_data = l1tol2net_io_managers_0_release_bits_data;
  assign L2BroadcastHub_1_io_inner_release_bits_client_id = l1tol2net_io_managers_0_release_bits_client_id;
  assign L2BroadcastHub_1_io_incoherent_0 = io_incoherent_0;
  assign L2BroadcastHub_1_io_outer_acquire_ready = ClientTileLinkEnqueuer_1_io_inner_acquire_ready;
  assign L2BroadcastHub_1_io_outer_probe_valid = ClientTileLinkEnqueuer_1_io_inner_probe_valid;
  assign L2BroadcastHub_1_io_outer_probe_bits_addr_block = ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block;
  assign L2BroadcastHub_1_io_outer_probe_bits_p_type = ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type;
  assign L2BroadcastHub_1_io_outer_release_ready = ClientTileLinkEnqueuer_1_io_inner_release_ready;
  assign L2BroadcastHub_1_io_outer_grant_valid = ClientTileLinkEnqueuer_1_io_inner_grant_valid;
  assign L2BroadcastHub_1_io_outer_grant_bits_addr_beat = ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  assign L2BroadcastHub_1_io_outer_grant_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  assign L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  assign L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type = ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  assign L2BroadcastHub_1_io_outer_grant_bits_g_type = ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  assign L2BroadcastHub_1_io_outer_grant_bits_data = ClientTileLinkEnqueuer_1_io_inner_grant_bits_data;
  assign L2BroadcastHub_1_io_outer_grant_bits_manager_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id;
  assign L2BroadcastHub_1_io_outer_finish_ready = ClientTileLinkEnqueuer_1_io_inner_finish_ready;
  assign mmioManager_clk = clk;
  assign mmioManager_reset = reset;
  assign mmioManager_io_inner_acquire_valid = l1tol2net_io_managers_1_acquire_valid;
  assign mmioManager_io_inner_acquire_bits_addr_block = l1tol2net_io_managers_1_acquire_bits_addr_block;
  assign mmioManager_io_inner_acquire_bits_client_xact_id = l1tol2net_io_managers_1_acquire_bits_client_xact_id;
  assign mmioManager_io_inner_acquire_bits_addr_beat = l1tol2net_io_managers_1_acquire_bits_addr_beat;
  assign mmioManager_io_inner_acquire_bits_is_builtin_type = l1tol2net_io_managers_1_acquire_bits_is_builtin_type;
  assign mmioManager_io_inner_acquire_bits_a_type = l1tol2net_io_managers_1_acquire_bits_a_type;
  assign mmioManager_io_inner_acquire_bits_union = l1tol2net_io_managers_1_acquire_bits_union;
  assign mmioManager_io_inner_acquire_bits_data = l1tol2net_io_managers_1_acquire_bits_data;
  assign mmioManager_io_inner_acquire_bits_client_id = l1tol2net_io_managers_1_acquire_bits_client_id;
  assign mmioManager_io_inner_grant_ready = l1tol2net_io_managers_1_grant_ready;
  assign mmioManager_io_inner_finish_valid = l1tol2net_io_managers_1_finish_valid;
  assign mmioManager_io_inner_finish_bits_manager_xact_id = l1tol2net_io_managers_1_finish_bits_manager_xact_id;
  assign mmioManager_io_inner_probe_ready = l1tol2net_io_managers_1_probe_ready;
  assign mmioManager_io_inner_release_valid = l1tol2net_io_managers_1_release_valid;
  assign mmioManager_io_inner_release_bits_addr_beat = l1tol2net_io_managers_1_release_bits_addr_beat;
  assign mmioManager_io_inner_release_bits_addr_block = l1tol2net_io_managers_1_release_bits_addr_block;
  assign mmioManager_io_inner_release_bits_client_xact_id = l1tol2net_io_managers_1_release_bits_client_xact_id;
  assign mmioManager_io_inner_release_bits_voluntary = l1tol2net_io_managers_1_release_bits_voluntary;
  assign mmioManager_io_inner_release_bits_r_type = l1tol2net_io_managers_1_release_bits_r_type;
  assign mmioManager_io_inner_release_bits_data = l1tol2net_io_managers_1_release_bits_data;
  assign mmioManager_io_inner_release_bits_client_id = l1tol2net_io_managers_1_release_bits_client_id;
  assign mmioManager_io_incoherent_0 = GEN_0;
  assign mmioManager_io_outer_acquire_ready = io_mmio_acquire_ready;
  assign mmioManager_io_outer_grant_valid = io_mmio_grant_valid;
  assign mmioManager_io_outer_grant_bits_addr_beat = io_mmio_grant_bits_addr_beat;
  assign mmioManager_io_outer_grant_bits_client_xact_id = io_mmio_grant_bits_client_xact_id;
  assign mmioManager_io_outer_grant_bits_manager_xact_id = io_mmio_grant_bits_manager_xact_id;
  assign mmioManager_io_outer_grant_bits_is_builtin_type = io_mmio_grant_bits_is_builtin_type;
  assign mmioManager_io_outer_grant_bits_g_type = io_mmio_grant_bits_g_type;
  assign mmioManager_io_outer_grant_bits_data = io_mmio_grant_bits_data;
  assign mem_ic_clk = clk;
  assign mem_ic_reset = reset;
  assign mem_ic_io_in_0_acquire_valid = ClientTileLinkIOUnwrapper_1_io_out_acquire_valid;
  assign mem_ic_io_in_0_acquire_bits_addr_block = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block;
  assign mem_ic_io_in_0_acquire_bits_client_xact_id = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id;
  assign mem_ic_io_in_0_acquire_bits_addr_beat = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat;
  assign mem_ic_io_in_0_acquire_bits_is_builtin_type = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type;
  assign mem_ic_io_in_0_acquire_bits_a_type = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type;
  assign mem_ic_io_in_0_acquire_bits_union = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union;
  assign mem_ic_io_in_0_acquire_bits_data = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data;
  assign mem_ic_io_in_0_grant_ready = ClientTileLinkIOUnwrapper_1_io_out_grant_ready;
  assign mem_ic_io_out_0_acquire_ready = NastiIOTileLinkIOConverter_1_io_tl_acquire_ready;
  assign mem_ic_io_out_0_grant_valid = NastiIOTileLinkIOConverter_1_io_tl_grant_valid;
  assign mem_ic_io_out_0_grant_bits_addr_beat = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat;
  assign mem_ic_io_out_0_grant_bits_client_xact_id = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id;
  assign mem_ic_io_out_0_grant_bits_manager_xact_id = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id;
  assign mem_ic_io_out_0_grant_bits_is_builtin_type = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type;
  assign mem_ic_io_out_0_grant_bits_g_type = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type;
  assign mem_ic_io_out_0_grant_bits_data = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data;
  assign ClientTileLinkIOUnwrapper_1_clk = clk;
  assign ClientTileLinkIOUnwrapper_1_reset = reset;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_valid = ClientTileLinkEnqueuer_1_io_outer_acquire_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  assign ClientTileLinkIOUnwrapper_1_io_in_probe_ready = ClientTileLinkEnqueuer_1_io_outer_probe_ready;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_valid = ClientTileLinkEnqueuer_1_io_outer_release_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat = ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block = ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary = ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type = ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_data = ClientTileLinkEnqueuer_1_io_outer_release_bits_data;
  assign ClientTileLinkIOUnwrapper_1_io_in_grant_ready = ClientTileLinkEnqueuer_1_io_outer_grant_ready;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_valid = ClientTileLinkEnqueuer_1_io_outer_finish_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id = ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id = ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_acquire_ready = mem_ic_io_in_0_acquire_ready;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_valid = mem_ic_io_in_0_grant_valid;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat = mem_ic_io_in_0_grant_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id = mem_ic_io_in_0_grant_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id = mem_ic_io_in_0_grant_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type = mem_ic_io_in_0_grant_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type = mem_ic_io_in_0_grant_bits_g_type;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data = mem_ic_io_in_0_grant_bits_data;
  assign ClientTileLinkEnqueuer_1_clk = clk;
  assign ClientTileLinkEnqueuer_1_reset = reset;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_valid = L2BroadcastHub_1_io_outer_acquire_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block = L2BroadcastHub_1_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id = L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat = L2BroadcastHub_1_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type = L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type = L2BroadcastHub_1_io_outer_acquire_bits_a_type;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union = L2BroadcastHub_1_io_outer_acquire_bits_union;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data = L2BroadcastHub_1_io_outer_acquire_bits_data;
  assign ClientTileLinkEnqueuer_1_io_inner_probe_ready = L2BroadcastHub_1_io_outer_probe_ready;
  assign ClientTileLinkEnqueuer_1_io_inner_release_valid = L2BroadcastHub_1_io_outer_release_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat = L2BroadcastHub_1_io_outer_release_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block = L2BroadcastHub_1_io_outer_release_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id = L2BroadcastHub_1_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary = L2BroadcastHub_1_io_outer_release_bits_voluntary;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type = L2BroadcastHub_1_io_outer_release_bits_r_type;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_data = L2BroadcastHub_1_io_outer_release_bits_data;
  assign ClientTileLinkEnqueuer_1_io_inner_grant_ready = L2BroadcastHub_1_io_outer_grant_ready;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_valid = L2BroadcastHub_1_io_outer_finish_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id = L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id = L2BroadcastHub_1_io_outer_finish_bits_manager_id;
  assign ClientTileLinkEnqueuer_1_io_outer_acquire_ready = ClientTileLinkIOUnwrapper_1_io_in_acquire_ready;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_valid = ClientTileLinkIOUnwrapper_1_io_in_probe_valid;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block = ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type = ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type;
  assign ClientTileLinkEnqueuer_1_io_outer_release_ready = ClientTileLinkIOUnwrapper_1_io_in_release_ready;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_valid = ClientTileLinkIOUnwrapper_1_io_in_grant_valid;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_data = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id;
  assign ClientTileLinkEnqueuer_1_io_outer_finish_ready = ClientTileLinkIOUnwrapper_1_io_in_finish_ready;
  assign NastiIOTileLinkIOConverter_1_clk = clk;
  assign NastiIOTileLinkIOConverter_1_reset = reset;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_valid = mem_ic_io_out_0_acquire_valid;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block = mem_ic_io_out_0_acquire_bits_addr_block;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id = mem_ic_io_out_0_acquire_bits_client_xact_id;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat = mem_ic_io_out_0_acquire_bits_addr_beat;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type = mem_ic_io_out_0_acquire_bits_is_builtin_type;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type = mem_ic_io_out_0_acquire_bits_a_type;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union = mem_ic_io_out_0_acquire_bits_union;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data = mem_ic_io_out_0_acquire_bits_data;
  assign NastiIOTileLinkIOConverter_1_io_tl_grant_ready = mem_ic_io_out_0_grant_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_aw_ready = Queue_16_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_w_ready = Queue_17_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_valid = Queue_19_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp = Queue_19_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id = Queue_19_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user = Queue_19_1_io_deq_bits_user;
  assign NastiIOTileLinkIOConverter_1_io_nasti_ar_ready = Queue_15_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_valid = Queue_18_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp = Queue_18_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data = Queue_18_1_io_deq_bits_data;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last = Queue_18_1_io_deq_bits_last;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id = Queue_18_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user = Queue_18_1_io_deq_bits_user;
  assign Queue_15_1_clk = clk;
  assign Queue_15_1_reset = reset;
  assign Queue_15_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_ar_valid;
  assign Queue_15_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr;
  assign Queue_15_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len;
  assign Queue_15_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size;
  assign Queue_15_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst;
  assign Queue_15_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock;
  assign Queue_15_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache;
  assign Queue_15_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot;
  assign Queue_15_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos;
  assign Queue_15_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region;
  assign Queue_15_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id;
  assign Queue_15_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user;
  assign Queue_15_1_io_deq_ready = io_mem_axi_0_ar_ready;
  assign Queue_16_1_clk = clk;
  assign Queue_16_1_reset = reset;
  assign Queue_16_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_aw_valid;
  assign Queue_16_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr;
  assign Queue_16_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len;
  assign Queue_16_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size;
  assign Queue_16_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst;
  assign Queue_16_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock;
  assign Queue_16_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache;
  assign Queue_16_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot;
  assign Queue_16_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos;
  assign Queue_16_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region;
  assign Queue_16_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id;
  assign Queue_16_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user;
  assign Queue_16_1_io_deq_ready = io_mem_axi_0_aw_ready;
  assign Queue_17_1_clk = clk;
  assign Queue_17_1_reset = reset;
  assign Queue_17_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_w_valid;
  assign Queue_17_1_io_enq_bits_data = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data;
  assign Queue_17_1_io_enq_bits_last = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last;
  assign Queue_17_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id;
  assign Queue_17_1_io_enq_bits_strb = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb;
  assign Queue_17_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user;
  assign Queue_17_1_io_deq_ready = io_mem_axi_0_w_ready;
  assign Queue_18_1_clk = clk;
  assign Queue_18_1_reset = reset;
  assign Queue_18_1_io_enq_valid = io_mem_axi_0_r_valid;
  assign Queue_18_1_io_enq_bits_resp = io_mem_axi_0_r_bits_resp;
  assign Queue_18_1_io_enq_bits_data = io_mem_axi_0_r_bits_data;
  assign Queue_18_1_io_enq_bits_last = io_mem_axi_0_r_bits_last;
  assign Queue_18_1_io_enq_bits_id = io_mem_axi_0_r_bits_id;
  assign Queue_18_1_io_enq_bits_user = io_mem_axi_0_r_bits_user;
  assign Queue_18_1_io_deq_ready = NastiIOTileLinkIOConverter_1_io_nasti_r_ready;
  assign Queue_19_1_clk = clk;
  assign Queue_19_1_reset = reset;
  assign Queue_19_1_io_enq_valid = io_mem_axi_0_b_valid;
  assign Queue_19_1_io_enq_bits_resp = io_mem_axi_0_b_bits_resp;
  assign Queue_19_1_io_enq_bits_id = io_mem_axi_0_b_bits_id;
  assign Queue_19_1_io_enq_bits_user = io_mem_axi_0_b_bits_user;
  assign Queue_19_1_io_deq_ready = NastiIOTileLinkIOConverter_1_io_nasti_b_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_1 = {1{$random}};
  GEN_0 = GEN_1[0:0];
  end
`endif
endmodule
module LockingRRArbiter_10(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_7;
  wire [2:0] GEN_1;
  wire [2:0] GEN_8;
  wire [1:0] GEN_2;
  wire [1:0] GEN_9;
  wire  GEN_3;
  wire  GEN_10;
  wire  GEN_4;
  wire  GEN_11;
  wire [3:0] GEN_5;
  wire [3:0] GEN_12;
  wire [63:0] GEN_6;
  wire [63:0] GEN_13;
  reg [2:0] T_610;
  reg [31:0] GEN_24;
  reg  T_612;
  reg [31:0] GEN_25;
  wire [2:0] GEN_20;
  wire  T_614;
  wire [2:0] T_622_0;
  wire [3:0] GEN_21;
  wire  T_624;
  wire  T_632_0;
  wire [3:0] GEN_22;
  wire  T_634;
  wire  T_637;
  wire  T_639;
  wire  T_640;
  wire [2:0] GEN_23;
  wire [3:0] T_644;
  wire [2:0] T_645;
  wire  GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  reg  lastGrant;
  reg [31:0] GEN_26;
  wire  GEN_17;
  wire  T_650;
  wire  T_652;
  wire  T_655;
  wire  T_659;
  wire  T_661;
  wire  T_665;
  wire  T_667;
  wire  T_668;
  wire  T_669;
  wire  T_672;
  wire  T_673;
  wire  GEN_18;
  wire  GEN_19;
  assign io_in_0_ready = T_669;
  assign io_in_1_ready = T_673;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_16;
  assign choice = GEN_19;
  assign GEN_0 = GEN_7;
  assign GEN_7 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_2 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_3 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_4 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_5 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_6 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_20 = {{2'd0}, 1'h0};
  assign T_614 = T_610 != GEN_20;
  assign T_622_0 = 3'h5;
  assign GEN_21 = {{1'd0}, T_622_0};
  assign T_624 = GEN_21 == io_out_bits_g_type;
  assign T_632_0 = 1'h0;
  assign GEN_22 = {{3'd0}, T_632_0};
  assign T_634 = GEN_22 == io_out_bits_g_type;
  assign T_637 = io_out_bits_is_builtin_type ? T_624 : T_634;
  assign T_639 = io_out_ready & io_out_valid;
  assign T_640 = T_639 & T_637;
  assign GEN_23 = {{2'd0}, 1'h1};
  assign T_644 = T_610 + GEN_23;
  assign T_645 = T_644[2:0];
  assign GEN_14 = T_640 ? io_chosen : T_612;
  assign GEN_15 = T_640 ? T_645 : T_610;
  assign GEN_16 = T_614 ? T_612 : choice;
  assign GEN_17 = T_639 ? io_chosen : lastGrant;
  assign T_650 = 1'h1 > lastGrant;
  assign T_652 = io_in_1_valid & T_650;
  assign T_655 = T_652 | io_in_0_valid;
  assign T_659 = T_652 == 1'h0;
  assign T_661 = T_655 == 1'h0;
  assign T_665 = T_650 | T_661;
  assign T_667 = T_612 == 1'h0;
  assign T_668 = T_614 ? T_667 : T_659;
  assign T_669 = T_668 & io_out_ready;
  assign T_672 = T_614 ? T_612 : T_665;
  assign T_673 = T_672 & io_out_ready;
  assign GEN_18 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_19 = T_652 ? 1'h1 : GEN_18;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_24 = {1{$random}};
  T_610 = GEN_24[2:0];
  GEN_25 = {1{$random}};
  T_612 = GEN_25[0:0];
  GEN_26 = {1{$random}};
  lastGrant = GEN_26[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_610 <= 3'h0;
    end else begin
      if(T_640) begin
        T_610 <= T_645;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_640) begin
        T_612 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_639) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIORouter(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data
);
  wire [2:0] T_1442;
  wire [28:0] T_1443;
  wire [31:0] T_1444;
  wire [31:0] GEN_2;
  wire  T_1448;
  wire [31:0] GEN_3;
  wire  T_1451;
  wire  T_1453;
  wire  T_1454;
  wire [1:0] acq_route;
  wire  T_1456;
  wire  T_1457;
  wire  GEN_0;
  wire  T_1459;
  wire  T_1460;
  wire  GEN_1;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_chosen;
  wire  T_1485;
  wire [1:0] GEN_4;
  wire  T_1487;
  wire  T_1488;
  wire  T_1489;
  wire  T_1491;
  LockingRRArbiter_10 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_1;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_1457;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign io_out_1_acquire_valid = T_1460;
  assign io_out_1_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_1_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_1_grant_ready = gnt_arb_io_in_1_ready;
  assign T_1442 = io_in_acquire_bits_union[11:9];
  assign T_1443 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_1444 = {T_1443,T_1442};
  assign GEN_2 = {{1'd0}, 31'h48000000};
  assign T_1448 = T_1444 < GEN_2;
  assign GEN_3 = {{1'd0}, 31'h60000000};
  assign T_1451 = GEN_3 <= T_1444;
  assign T_1453 = T_1444 < 32'h80000000;
  assign T_1454 = T_1451 & T_1453;
  assign acq_route = {T_1454,T_1448};
  assign T_1456 = acq_route[0];
  assign T_1457 = io_in_acquire_valid & T_1456;
  assign GEN_0 = T_1456 ? io_out_0_acquire_ready : 1'h0;
  assign T_1459 = acq_route[1];
  assign T_1460 = io_in_acquire_valid & T_1459;
  assign GEN_1 = T_1459 ? io_out_1_acquire_ready : GEN_0;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_in_1_valid = io_out_1_grant_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = io_out_1_grant_bits_g_type;
  assign gnt_arb_io_in_1_bits_data = io_out_1_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_1485 = io_in_acquire_valid == 1'h0;
  assign GEN_4 = {{1'd0}, 1'h0};
  assign T_1487 = acq_route != GEN_4;
  assign T_1488 = T_1485 | T_1487;
  assign T_1489 = T_1488 | reset;
  assign T_1491 = T_1489 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1491) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at Interconnect.scala:219 assert(!io.in.acquire.valid || acq_route.orR, \"No valid route\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1491) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1491) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_1_clk;
  wire  ClientUncachedTileLinkIORouter_1_reset;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_data;
  ClientUncachedTileLinkIORouter ClientUncachedTileLinkIORouter_1 (
    .clk(ClientUncachedTileLinkIORouter_1_clk),
    .reset(ClientUncachedTileLinkIORouter_1_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_1_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(ClientUncachedTileLinkIORouter_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(ClientUncachedTileLinkIORouter_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_1_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_1_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = ClientUncachedTileLinkIORouter_1_io_out_1_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_clk = clk;
  assign ClientUncachedTileLinkIORouter_1_reset = reset;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_1_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
endmodule
module LockingRRArbiter_11(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [1:0] io_in_2_bits_client_xact_id,
  input   io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [1:0] io_in_3_bits_client_xact_id,
  input   io_in_3_bits_manager_xact_id,
  input   io_in_3_bits_is_builtin_type,
  input  [3:0] io_in_3_bits_g_type,
  input  [63:0] io_in_3_bits_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_addr_beat,
  input  [1:0] io_in_4_bits_client_xact_id,
  input   io_in_4_bits_manager_xact_id,
  input   io_in_4_bits_is_builtin_type,
  input  [3:0] io_in_4_bits_g_type,
  input  [63:0] io_in_4_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_47;
  wire  GEN_7;
  wire [2:0] GEN_48;
  wire  GEN_8;
  wire [2:0] GEN_49;
  wire  GEN_9;
  wire  GEN_10;
  wire [2:0] GEN_1;
  wire [2:0] GEN_11;
  wire [2:0] GEN_12;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [1:0] GEN_2;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire  GEN_3;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_4;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire [3:0] GEN_5;
  wire [3:0] GEN_27;
  wire [3:0] GEN_28;
  wire [3:0] GEN_29;
  wire [3:0] GEN_30;
  wire [63:0] GEN_6;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  reg [2:0] T_886;
  reg [31:0] GEN_50;
  reg [2:0] T_888;
  reg [31:0] GEN_51;
  wire [2:0] GEN_68;
  wire  T_890;
  wire [2:0] T_898_0;
  wire [3:0] GEN_69;
  wire  T_900;
  wire  T_908_0;
  wire [3:0] GEN_70;
  wire  T_910;
  wire  T_913;
  wire  T_915;
  wire  T_916;
  wire [3:0] T_920;
  wire [2:0] T_921;
  wire [2:0] GEN_35;
  wire [2:0] GEN_36;
  wire [2:0] GEN_37;
  reg [2:0] lastGrant;
  reg [31:0] GEN_52;
  wire [2:0] GEN_38;
  wire  T_926;
  wire  T_928;
  wire  T_930;
  wire  T_932;
  wire  T_934;
  wire  T_935;
  wire  T_936;
  wire  T_937;
  wire  T_940;
  wire  T_941;
  wire  T_942;
  wire  T_943;
  wire  T_944;
  wire  T_945;
  wire  T_946;
  wire  T_950;
  wire  T_952;
  wire  T_954;
  wire  T_956;
  wire  T_958;
  wire  T_960;
  wire  T_962;
  wire  T_964;
  wire  T_968;
  wire  T_969;
  wire  T_970;
  wire  T_971;
  wire  T_972;
  wire  T_973;
  wire  T_974;
  wire  T_976;
  wire  T_977;
  wire  T_978;
  wire  T_980;
  wire  T_981;
  wire  T_982;
  wire  T_984;
  wire  T_985;
  wire  T_986;
  wire  T_988;
  wire  T_989;
  wire  T_990;
  wire  T_992;
  wire  T_993;
  wire  T_994;
  wire [2:0] GEN_39;
  wire [2:0] GEN_40;
  wire [2:0] GEN_41;
  wire [2:0] GEN_42;
  wire [2:0] GEN_43;
  wire [2:0] GEN_44;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  assign io_in_0_ready = T_978;
  assign io_in_1_ready = T_982;
  assign io_in_2_ready = T_986;
  assign io_in_3_ready = T_990;
  assign io_in_4_ready = T_994;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_37;
  assign choice = GEN_46;
  assign GEN_0 = GEN_10;
  assign GEN_47 = {{2'd0}, 1'h1};
  assign GEN_7 = GEN_47 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_48 = {{1'd0}, 2'h2};
  assign GEN_8 = GEN_48 == io_chosen ? io_in_2_valid : GEN_7;
  assign GEN_49 = {{1'd0}, 2'h3};
  assign GEN_9 = GEN_49 == io_chosen ? io_in_3_valid : GEN_8;
  assign GEN_10 = 3'h4 == io_chosen ? io_in_4_valid : GEN_9;
  assign GEN_1 = GEN_14;
  assign GEN_11 = GEN_47 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_12 = GEN_48 == io_chosen ? io_in_2_bits_addr_beat : GEN_11;
  assign GEN_13 = GEN_49 == io_chosen ? io_in_3_bits_addr_beat : GEN_12;
  assign GEN_14 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_13;
  assign GEN_2 = GEN_18;
  assign GEN_15 = GEN_47 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_16 = GEN_48 == io_chosen ? io_in_2_bits_client_xact_id : GEN_15;
  assign GEN_17 = GEN_49 == io_chosen ? io_in_3_bits_client_xact_id : GEN_16;
  assign GEN_18 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_17;
  assign GEN_3 = GEN_22;
  assign GEN_19 = GEN_47 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_20 = GEN_48 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_19;
  assign GEN_21 = GEN_49 == io_chosen ? io_in_3_bits_manager_xact_id : GEN_20;
  assign GEN_22 = 3'h4 == io_chosen ? io_in_4_bits_manager_xact_id : GEN_21;
  assign GEN_4 = GEN_26;
  assign GEN_23 = GEN_47 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_24 = GEN_48 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_23;
  assign GEN_25 = GEN_49 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_24;
  assign GEN_26 = 3'h4 == io_chosen ? io_in_4_bits_is_builtin_type : GEN_25;
  assign GEN_5 = GEN_30;
  assign GEN_27 = GEN_47 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_28 = GEN_48 == io_chosen ? io_in_2_bits_g_type : GEN_27;
  assign GEN_29 = GEN_49 == io_chosen ? io_in_3_bits_g_type : GEN_28;
  assign GEN_30 = 3'h4 == io_chosen ? io_in_4_bits_g_type : GEN_29;
  assign GEN_6 = GEN_34;
  assign GEN_31 = GEN_47 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_32 = GEN_48 == io_chosen ? io_in_2_bits_data : GEN_31;
  assign GEN_33 = GEN_49 == io_chosen ? io_in_3_bits_data : GEN_32;
  assign GEN_34 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_33;
  assign GEN_68 = {{2'd0}, 1'h0};
  assign T_890 = T_886 != GEN_68;
  assign T_898_0 = 3'h5;
  assign GEN_69 = {{1'd0}, T_898_0};
  assign T_900 = GEN_69 == io_out_bits_g_type;
  assign T_908_0 = 1'h0;
  assign GEN_70 = {{3'd0}, T_908_0};
  assign T_910 = GEN_70 == io_out_bits_g_type;
  assign T_913 = io_out_bits_is_builtin_type ? T_900 : T_910;
  assign T_915 = io_out_ready & io_out_valid;
  assign T_916 = T_915 & T_913;
  assign T_920 = T_886 + GEN_47;
  assign T_921 = T_920[2:0];
  assign GEN_35 = T_916 ? io_chosen : T_888;
  assign GEN_36 = T_916 ? T_921 : T_886;
  assign GEN_37 = T_890 ? T_888 : choice;
  assign GEN_38 = T_915 ? io_chosen : lastGrant;
  assign T_926 = GEN_47 > lastGrant;
  assign T_928 = GEN_48 > lastGrant;
  assign T_930 = GEN_49 > lastGrant;
  assign T_932 = 3'h4 > lastGrant;
  assign T_934 = io_in_1_valid & T_926;
  assign T_935 = io_in_2_valid & T_928;
  assign T_936 = io_in_3_valid & T_930;
  assign T_937 = io_in_4_valid & T_932;
  assign T_940 = T_934 | T_935;
  assign T_941 = T_940 | T_936;
  assign T_942 = T_941 | T_937;
  assign T_943 = T_942 | io_in_0_valid;
  assign T_944 = T_943 | io_in_1_valid;
  assign T_945 = T_944 | io_in_2_valid;
  assign T_946 = T_945 | io_in_3_valid;
  assign T_950 = T_934 == 1'h0;
  assign T_952 = T_940 == 1'h0;
  assign T_954 = T_941 == 1'h0;
  assign T_956 = T_942 == 1'h0;
  assign T_958 = T_943 == 1'h0;
  assign T_960 = T_944 == 1'h0;
  assign T_962 = T_945 == 1'h0;
  assign T_964 = T_946 == 1'h0;
  assign T_968 = T_926 | T_958;
  assign T_969 = T_950 & T_928;
  assign T_970 = T_969 | T_960;
  assign T_971 = T_952 & T_930;
  assign T_972 = T_971 | T_962;
  assign T_973 = T_954 & T_932;
  assign T_974 = T_973 | T_964;
  assign T_976 = T_888 == GEN_68;
  assign T_977 = T_890 ? T_976 : T_956;
  assign T_978 = T_977 & io_out_ready;
  assign T_980 = T_888 == GEN_47;
  assign T_981 = T_890 ? T_980 : T_968;
  assign T_982 = T_981 & io_out_ready;
  assign T_984 = T_888 == GEN_48;
  assign T_985 = T_890 ? T_984 : T_970;
  assign T_986 = T_985 & io_out_ready;
  assign T_988 = T_888 == GEN_49;
  assign T_989 = T_890 ? T_988 : T_972;
  assign T_990 = T_989 & io_out_ready;
  assign T_992 = T_888 == 3'h4;
  assign T_993 = T_890 ? T_992 : T_974;
  assign T_994 = T_993 & io_out_ready;
  assign GEN_39 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_40 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_39;
  assign GEN_41 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_40;
  assign GEN_42 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_41;
  assign GEN_43 = T_937 ? 3'h4 : GEN_42;
  assign GEN_44 = T_936 ? {{1'd0}, 2'h3} : GEN_43;
  assign GEN_45 = T_935 ? {{1'd0}, 2'h2} : GEN_44;
  assign GEN_46 = T_934 ? {{2'd0}, 1'h1} : GEN_45;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_50 = {1{$random}};
  T_886 = GEN_50[2:0];
  GEN_51 = {1{$random}};
  T_888 = GEN_51[2:0];
  GEN_52 = {1{$random}};
  lastGrant = GEN_52[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_886 <= 3'h0;
    end else begin
      if(T_916) begin
        T_886 <= T_921;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_916) begin
        T_888 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_915) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIORouter_1(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data
);
  wire [2:0] T_2051;
  wire [28:0] T_2052;
  wire [31:0] T_2053;
  wire [31:0] GEN_5;
  wire  T_2057;
  wire  T_2060;
  wire [31:0] GEN_7;
  wire  T_2062;
  wire  T_2063;
  wire  T_2065;
  wire [31:0] GEN_9;
  wire  T_2067;
  wire  T_2068;
  wire [31:0] GEN_10;
  wire  T_2070;
  wire [31:0] GEN_11;
  wire  T_2072;
  wire  T_2073;
  wire  T_2075;
  wire [31:0] GEN_13;
  wire  T_2077;
  wire  T_2078;
  wire [1:0] T_2079;
  wire [1:0] T_2080;
  wire [2:0] T_2081;
  wire [4:0] acq_route;
  wire  T_2083;
  wire  T_2084;
  wire  GEN_0;
  wire  T_2086;
  wire  T_2087;
  wire  GEN_1;
  wire  T_2089;
  wire  T_2090;
  wire  GEN_2;
  wire  T_2092;
  wire  T_2093;
  wire  GEN_3;
  wire  T_2095;
  wire  T_2096;
  wire  GEN_4;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_2_ready;
  wire  gnt_arb_io_in_2_valid;
  wire [2:0] gnt_arb_io_in_2_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_2_bits_client_xact_id;
  wire  gnt_arb_io_in_2_bits_manager_xact_id;
  wire  gnt_arb_io_in_2_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_2_bits_g_type;
  wire [63:0] gnt_arb_io_in_2_bits_data;
  wire  gnt_arb_io_in_3_ready;
  wire  gnt_arb_io_in_3_valid;
  wire [2:0] gnt_arb_io_in_3_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_3_bits_client_xact_id;
  wire  gnt_arb_io_in_3_bits_manager_xact_id;
  wire  gnt_arb_io_in_3_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_3_bits_g_type;
  wire [63:0] gnt_arb_io_in_3_bits_data;
  wire  gnt_arb_io_in_4_ready;
  wire  gnt_arb_io_in_4_valid;
  wire [2:0] gnt_arb_io_in_4_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_4_bits_client_xact_id;
  wire  gnt_arb_io_in_4_bits_manager_xact_id;
  wire  gnt_arb_io_in_4_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_4_bits_g_type;
  wire [63:0] gnt_arb_io_in_4_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire [2:0] gnt_arb_io_chosen;
  wire  T_2121;
  wire [4:0] GEN_14;
  wire  T_2123;
  wire  T_2124;
  wire  T_2125;
  wire  T_2127;
  LockingRRArbiter_11 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_2_ready(gnt_arb_io_in_2_ready),
    .io_in_2_valid(gnt_arb_io_in_2_valid),
    .io_in_2_bits_addr_beat(gnt_arb_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(gnt_arb_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(gnt_arb_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(gnt_arb_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(gnt_arb_io_in_2_bits_g_type),
    .io_in_2_bits_data(gnt_arb_io_in_2_bits_data),
    .io_in_3_ready(gnt_arb_io_in_3_ready),
    .io_in_3_valid(gnt_arb_io_in_3_valid),
    .io_in_3_bits_addr_beat(gnt_arb_io_in_3_bits_addr_beat),
    .io_in_3_bits_client_xact_id(gnt_arb_io_in_3_bits_client_xact_id),
    .io_in_3_bits_manager_xact_id(gnt_arb_io_in_3_bits_manager_xact_id),
    .io_in_3_bits_is_builtin_type(gnt_arb_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_g_type(gnt_arb_io_in_3_bits_g_type),
    .io_in_3_bits_data(gnt_arb_io_in_3_bits_data),
    .io_in_4_ready(gnt_arb_io_in_4_ready),
    .io_in_4_valid(gnt_arb_io_in_4_valid),
    .io_in_4_bits_addr_beat(gnt_arb_io_in_4_bits_addr_beat),
    .io_in_4_bits_client_xact_id(gnt_arb_io_in_4_bits_client_xact_id),
    .io_in_4_bits_manager_xact_id(gnt_arb_io_in_4_bits_manager_xact_id),
    .io_in_4_bits_is_builtin_type(gnt_arb_io_in_4_bits_is_builtin_type),
    .io_in_4_bits_g_type(gnt_arb_io_in_4_bits_g_type),
    .io_in_4_bits_data(gnt_arb_io_in_4_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_4;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_2084;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign io_out_1_acquire_valid = T_2087;
  assign io_out_1_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_1_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_1_grant_ready = gnt_arb_io_in_1_ready;
  assign io_out_2_acquire_valid = T_2090;
  assign io_out_2_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_2_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_2_grant_ready = gnt_arb_io_in_2_ready;
  assign io_out_3_acquire_valid = T_2093;
  assign io_out_3_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_3_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_3_grant_ready = gnt_arb_io_in_3_ready;
  assign io_out_4_acquire_valid = T_2096;
  assign io_out_4_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_4_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_4_grant_ready = gnt_arb_io_in_4_ready;
  assign T_2051 = io_in_acquire_bits_union[11:9];
  assign T_2052 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_2053 = {T_2052,T_2051};
  assign GEN_5 = {{19'd0}, 13'h1000};
  assign T_2057 = T_2053 < GEN_5;
  assign T_2060 = GEN_5 <= T_2053;
  assign GEN_7 = {{18'd0}, 14'h2000};
  assign T_2062 = T_2053 < GEN_7;
  assign T_2063 = T_2060 & T_2062;
  assign T_2065 = GEN_7 <= T_2053;
  assign GEN_9 = {{17'd0}, 15'h4000};
  assign T_2067 = T_2053 < GEN_9;
  assign T_2068 = T_2065 & T_2067;
  assign GEN_10 = {{1'd0}, 31'h40000000};
  assign T_2070 = GEN_10 <= T_2053;
  assign GEN_11 = {{1'd0}, 31'h44000000};
  assign T_2072 = T_2053 < GEN_11;
  assign T_2073 = T_2070 & T_2072;
  assign T_2075 = GEN_11 <= T_2053;
  assign GEN_13 = {{1'd0}, 31'h48000000};
  assign T_2077 = T_2053 < GEN_13;
  assign T_2078 = T_2075 & T_2077;
  assign T_2079 = {T_2063,T_2057};
  assign T_2080 = {T_2078,T_2073};
  assign T_2081 = {T_2080,T_2068};
  assign acq_route = {T_2081,T_2079};
  assign T_2083 = acq_route[0];
  assign T_2084 = io_in_acquire_valid & T_2083;
  assign GEN_0 = T_2083 ? io_out_0_acquire_ready : 1'h0;
  assign T_2086 = acq_route[1];
  assign T_2087 = io_in_acquire_valid & T_2086;
  assign GEN_1 = T_2086 ? io_out_1_acquire_ready : GEN_0;
  assign T_2089 = acq_route[2];
  assign T_2090 = io_in_acquire_valid & T_2089;
  assign GEN_2 = T_2089 ? io_out_2_acquire_ready : GEN_1;
  assign T_2092 = acq_route[3];
  assign T_2093 = io_in_acquire_valid & T_2092;
  assign GEN_3 = T_2092 ? io_out_3_acquire_ready : GEN_2;
  assign T_2095 = acq_route[4];
  assign T_2096 = io_in_acquire_valid & T_2095;
  assign GEN_4 = T_2095 ? io_out_4_acquire_ready : GEN_3;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_in_1_valid = io_out_1_grant_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = io_out_1_grant_bits_g_type;
  assign gnt_arb_io_in_1_bits_data = io_out_1_grant_bits_data;
  assign gnt_arb_io_in_2_valid = io_out_2_grant_valid;
  assign gnt_arb_io_in_2_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign gnt_arb_io_in_2_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign gnt_arb_io_in_2_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_2_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_2_bits_g_type = io_out_2_grant_bits_g_type;
  assign gnt_arb_io_in_2_bits_data = io_out_2_grant_bits_data;
  assign gnt_arb_io_in_3_valid = io_out_3_grant_valid;
  assign gnt_arb_io_in_3_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign gnt_arb_io_in_3_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign gnt_arb_io_in_3_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_3_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_3_bits_g_type = io_out_3_grant_bits_g_type;
  assign gnt_arb_io_in_3_bits_data = io_out_3_grant_bits_data;
  assign gnt_arb_io_in_4_valid = io_out_4_grant_valid;
  assign gnt_arb_io_in_4_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign gnt_arb_io_in_4_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign gnt_arb_io_in_4_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_4_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_4_bits_g_type = io_out_4_grant_bits_g_type;
  assign gnt_arb_io_in_4_bits_data = io_out_4_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_2121 = io_in_acquire_valid == 1'h0;
  assign GEN_14 = {{4'd0}, 1'h0};
  assign T_2123 = acq_route != GEN_14;
  assign T_2124 = T_2121 | T_2123;
  assign T_2125 = T_2124 | reset;
  assign T_2127 = T_2125 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2127) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at Interconnect.scala:219 assert(!io.in.acquire.valid || acq_route.orR, \"No valid route\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2127) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_2127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_1_1_clk;
  wire  ClientUncachedTileLinkIORouter_1_1_reset;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_data;
  ClientUncachedTileLinkIORouter_1 ClientUncachedTileLinkIORouter_1_1 (
    .clk(ClientUncachedTileLinkIORouter_1_1_clk),
    .reset(ClientUncachedTileLinkIORouter_1_1_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready),
    .io_out_2_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready),
    .io_out_3_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_ready),
    .io_out_4_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready;
  assign io_out_4_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_valid;
  assign io_out_4_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_union;
  assign io_out_4_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_bits_data;
  assign io_out_4_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_1_clk = clk;
  assign ClientUncachedTileLinkIORouter_1_1_reset = reset;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid = io_out_2_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid = io_out_3_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_4_acquire_ready = io_out_4_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_valid = io_out_4_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_g_type = io_out_4_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_4_grant_bits_data = io_out_4_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [11:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [11:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  xbar_io_out_1_acquire_ready;
  wire  xbar_io_out_1_acquire_valid;
  wire [25:0] xbar_io_out_1_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_1_acquire_bits_addr_beat;
  wire  xbar_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_1_acquire_bits_a_type;
  wire [11:0] xbar_io_out_1_acquire_bits_union;
  wire [63:0] xbar_io_out_1_acquire_bits_data;
  wire  xbar_io_out_1_grant_ready;
  wire  xbar_io_out_1_grant_valid;
  wire [2:0] xbar_io_out_1_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_1_grant_bits_client_xact_id;
  wire  xbar_io_out_1_grant_bits_manager_xact_id;
  wire  xbar_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_1_grant_bits_g_type;
  wire [63:0] xbar_io_out_1_grant_bits_data;
  wire  xbar_io_out_2_acquire_ready;
  wire  xbar_io_out_2_acquire_valid;
  wire [25:0] xbar_io_out_2_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_2_acquire_bits_addr_beat;
  wire  xbar_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_2_acquire_bits_a_type;
  wire [11:0] xbar_io_out_2_acquire_bits_union;
  wire [63:0] xbar_io_out_2_acquire_bits_data;
  wire  xbar_io_out_2_grant_ready;
  wire  xbar_io_out_2_grant_valid;
  wire [2:0] xbar_io_out_2_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_2_grant_bits_client_xact_id;
  wire  xbar_io_out_2_grant_bits_manager_xact_id;
  wire  xbar_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_2_grant_bits_g_type;
  wire [63:0] xbar_io_out_2_grant_bits_data;
  wire  xbar_io_out_3_acquire_ready;
  wire  xbar_io_out_3_acquire_valid;
  wire [25:0] xbar_io_out_3_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_3_acquire_bits_addr_beat;
  wire  xbar_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_3_acquire_bits_a_type;
  wire [11:0] xbar_io_out_3_acquire_bits_union;
  wire [63:0] xbar_io_out_3_acquire_bits_data;
  wire  xbar_io_out_3_grant_ready;
  wire  xbar_io_out_3_grant_valid;
  wire [2:0] xbar_io_out_3_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_3_grant_bits_client_xact_id;
  wire  xbar_io_out_3_grant_bits_manager_xact_id;
  wire  xbar_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_3_grant_bits_g_type;
  wire [63:0] xbar_io_out_3_grant_bits_data;
  wire  xbar_io_out_4_acquire_ready;
  wire  xbar_io_out_4_acquire_valid;
  wire [25:0] xbar_io_out_4_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_4_acquire_bits_addr_beat;
  wire  xbar_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_4_acquire_bits_a_type;
  wire [11:0] xbar_io_out_4_acquire_bits_union;
  wire [63:0] xbar_io_out_4_acquire_bits_data;
  wire  xbar_io_out_4_grant_ready;
  wire  xbar_io_out_4_grant_valid;
  wire [2:0] xbar_io_out_4_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_4_grant_bits_client_xact_id;
  wire  xbar_io_out_4_grant_bits_manager_xact_id;
  wire  xbar_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_4_grant_bits_g_type;
  wire [63:0] xbar_io_out_4_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar_1 xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(xbar_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(xbar_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(xbar_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(xbar_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(xbar_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(xbar_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(xbar_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(xbar_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(xbar_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(xbar_io_out_1_grant_ready),
    .io_out_1_grant_valid(xbar_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(xbar_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(xbar_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(xbar_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(xbar_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(xbar_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(xbar_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(xbar_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(xbar_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(xbar_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(xbar_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(xbar_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(xbar_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(xbar_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(xbar_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(xbar_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(xbar_io_out_2_grant_ready),
    .io_out_2_grant_valid(xbar_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(xbar_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(xbar_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(xbar_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(xbar_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(xbar_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(xbar_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(xbar_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(xbar_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(xbar_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(xbar_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(xbar_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(xbar_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(xbar_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(xbar_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(xbar_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(xbar_io_out_3_grant_ready),
    .io_out_3_grant_valid(xbar_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(xbar_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(xbar_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(xbar_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(xbar_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(xbar_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(xbar_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(xbar_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(xbar_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(xbar_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(xbar_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(xbar_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(xbar_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(xbar_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(xbar_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(xbar_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(xbar_io_out_4_grant_ready),
    .io_out_4_grant_valid(xbar_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(xbar_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(xbar_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(xbar_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(xbar_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(xbar_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(xbar_io_out_4_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = xbar_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = xbar_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = xbar_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = xbar_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = xbar_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = xbar_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = xbar_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = xbar_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = xbar_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = xbar_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = xbar_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = xbar_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = xbar_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = xbar_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = xbar_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = xbar_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = xbar_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = xbar_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = xbar_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = xbar_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = xbar_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = xbar_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = xbar_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = xbar_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = xbar_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = xbar_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = xbar_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = xbar_io_out_3_grant_ready;
  assign io_out_4_acquire_valid = xbar_io_out_4_acquire_valid;
  assign io_out_4_acquire_bits_addr_block = xbar_io_out_4_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = xbar_io_out_4_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = xbar_io_out_4_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = xbar_io_out_4_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = xbar_io_out_4_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = xbar_io_out_4_acquire_bits_union;
  assign io_out_4_acquire_bits_data = xbar_io_out_4_acquire_bits_data;
  assign io_out_4_grant_ready = xbar_io_out_4_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = io_out_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign xbar_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign xbar_io_out_1_grant_valid = io_out_1_grant_valid;
  assign xbar_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign xbar_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign xbar_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign xbar_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign xbar_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign xbar_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign xbar_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign xbar_io_out_2_grant_valid = io_out_2_grant_valid;
  assign xbar_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign xbar_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign xbar_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign xbar_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign xbar_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign xbar_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign xbar_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign xbar_io_out_3_grant_valid = io_out_3_grant_valid;
  assign xbar_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign xbar_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign xbar_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign xbar_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign xbar_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign xbar_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
  assign xbar_io_out_4_acquire_ready = io_out_4_acquire_ready;
  assign xbar_io_out_4_grant_valid = io_out_4_grant_valid;
  assign xbar_io_out_4_grant_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign xbar_io_out_4_grant_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign xbar_io_out_4_grant_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign xbar_io_out_4_grant_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign xbar_io_out_4_grant_bits_g_type = io_out_4_grant_bits_g_type;
  assign xbar_io_out_4_grant_bits_data = io_out_4_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data,
  input   io_out_5_acquire_ready,
  output  io_out_5_acquire_valid,
  output [25:0] io_out_5_acquire_bits_addr_block,
  output [1:0] io_out_5_acquire_bits_client_xact_id,
  output [2:0] io_out_5_acquire_bits_addr_beat,
  output  io_out_5_acquire_bits_is_builtin_type,
  output [2:0] io_out_5_acquire_bits_a_type,
  output [11:0] io_out_5_acquire_bits_union,
  output [63:0] io_out_5_acquire_bits_data,
  output  io_out_5_grant_ready,
  input   io_out_5_grant_valid,
  input  [2:0] io_out_5_grant_bits_addr_beat,
  input  [1:0] io_out_5_grant_bits_client_xact_id,
  input   io_out_5_grant_bits_manager_xact_id,
  input   io_out_5_grant_bits_is_builtin_type,
  input  [3:0] io_out_5_grant_bits_g_type,
  input  [63:0] io_out_5_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [11:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [11:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  xbar_io_out_1_acquire_ready;
  wire  xbar_io_out_1_acquire_valid;
  wire [25:0] xbar_io_out_1_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_1_acquire_bits_addr_beat;
  wire  xbar_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_1_acquire_bits_a_type;
  wire [11:0] xbar_io_out_1_acquire_bits_union;
  wire [63:0] xbar_io_out_1_acquire_bits_data;
  wire  xbar_io_out_1_grant_ready;
  wire  xbar_io_out_1_grant_valid;
  wire [2:0] xbar_io_out_1_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_1_grant_bits_client_xact_id;
  wire  xbar_io_out_1_grant_bits_manager_xact_id;
  wire  xbar_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_1_grant_bits_g_type;
  wire [63:0] xbar_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_clk;
  wire  TileLinkRecursiveInterconnect_1_1_reset;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_4_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_4_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(xbar_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(xbar_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(xbar_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(xbar_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(xbar_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(xbar_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(xbar_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(xbar_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(xbar_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(xbar_io_out_1_grant_ready),
    .io_out_1_grant_valid(xbar_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(xbar_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(xbar_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(xbar_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(xbar_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(xbar_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(xbar_io_out_1_grant_bits_data)
  );
  TileLinkRecursiveInterconnect_1 TileLinkRecursiveInterconnect_1_1 (
    .clk(TileLinkRecursiveInterconnect_1_1_clk),
    .reset(TileLinkRecursiveInterconnect_1_1_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_4_grant_ready),
    .io_out_4_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready;
  assign io_out_4_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_valid;
  assign io_out_4_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_union;
  assign io_out_4_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_bits_data;
  assign io_out_4_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_4_grant_ready;
  assign io_out_5_acquire_valid = xbar_io_out_1_acquire_valid;
  assign io_out_5_acquire_bits_addr_block = xbar_io_out_1_acquire_bits_addr_block;
  assign io_out_5_acquire_bits_client_xact_id = xbar_io_out_1_acquire_bits_client_xact_id;
  assign io_out_5_acquire_bits_addr_beat = xbar_io_out_1_acquire_bits_addr_beat;
  assign io_out_5_acquire_bits_is_builtin_type = xbar_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_5_acquire_bits_a_type = xbar_io_out_1_acquire_bits_a_type;
  assign io_out_5_acquire_bits_union = xbar_io_out_1_acquire_bits_union;
  assign io_out_5_acquire_bits_data = xbar_io_out_1_acquire_bits_data;
  assign io_out_5_grant_ready = xbar_io_out_1_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data;
  assign xbar_io_out_1_acquire_ready = io_out_5_acquire_ready;
  assign xbar_io_out_1_grant_valid = io_out_5_grant_valid;
  assign xbar_io_out_1_grant_bits_addr_beat = io_out_5_grant_bits_addr_beat;
  assign xbar_io_out_1_grant_bits_client_xact_id = io_out_5_grant_bits_client_xact_id;
  assign xbar_io_out_1_grant_bits_manager_xact_id = io_out_5_grant_bits_manager_xact_id;
  assign xbar_io_out_1_grant_bits_is_builtin_type = io_out_5_grant_bits_is_builtin_type;
  assign xbar_io_out_1_grant_bits_g_type = io_out_5_grant_bits_g_type;
  assign xbar_io_out_1_grant_bits_data = io_out_5_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_clk = clk;
  assign TileLinkRecursiveInterconnect_1_1_reset = reset;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready = xbar_io_out_0_grant_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid = io_out_2_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid = io_out_3_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_4_acquire_ready = io_out_4_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_4_grant_valid = io_out_4_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_g_type = io_out_4_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_4_grant_bits_data = io_out_4_grant_bits_data;
endmodule
module Queue_20(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [25:0] io_enq_bits_addr_block,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input  [11:0] io_enq_bits_union,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [25:0] io_deq_bits_addr_block,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [11:0] io_deq_bits_union,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [25:0] ram_addr_block [0:0];
  reg [31:0] GEN_0;
  wire [25:0] ram_addr_block_T_254_data;
  wire  ram_addr_block_T_254_addr;
  wire  ram_addr_block_T_254_en;
  wire [25:0] ram_addr_block_T_224_data;
  wire  ram_addr_block_T_224_addr;
  wire  ram_addr_block_T_224_mask;
  wire  ram_addr_block_T_224_en;
  reg [1:0] ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_client_xact_id_T_254_data;
  wire  ram_client_xact_id_T_254_addr;
  wire  ram_client_xact_id_T_254_en;
  wire [1:0] ram_client_xact_id_T_224_data;
  wire  ram_client_xact_id_T_224_addr;
  wire  ram_client_xact_id_T_224_mask;
  wire  ram_client_xact_id_T_224_en;
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_addr_beat_T_254_data;
  wire  ram_addr_beat_T_254_addr;
  wire  ram_addr_beat_T_254_en;
  wire [2:0] ram_addr_beat_T_224_data;
  wire  ram_addr_beat_T_224_addr;
  wire  ram_addr_beat_T_224_mask;
  wire  ram_addr_beat_T_224_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_254_data;
  wire  ram_is_builtin_type_T_254_addr;
  wire  ram_is_builtin_type_T_254_en;
  wire  ram_is_builtin_type_T_224_data;
  wire  ram_is_builtin_type_T_224_addr;
  wire  ram_is_builtin_type_T_224_mask;
  wire  ram_is_builtin_type_T_224_en;
  reg [2:0] ram_a_type [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_254_data;
  wire  ram_a_type_T_254_addr;
  wire  ram_a_type_T_254_en;
  wire [2:0] ram_a_type_T_224_data;
  wire  ram_a_type_T_224_addr;
  wire  ram_a_type_T_224_mask;
  wire  ram_a_type_T_224_en;
  reg [11:0] ram_union [0:0];
  reg [31:0] GEN_5;
  wire [11:0] ram_union_T_254_data;
  wire  ram_union_T_254_addr;
  wire  ram_union_T_254_en;
  wire [11:0] ram_union_T_224_data;
  wire  ram_union_T_224_addr;
  wire  ram_union_T_224_mask;
  wire  ram_union_T_224_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_6;
  wire [63:0] ram_data_T_254_data;
  wire  ram_data_T_254_addr;
  wire  ram_data_T_254_en;
  wire [63:0] ram_data_T_224_data;
  wire  ram_data_T_224_addr;
  wire  ram_data_T_224_mask;
  wire  ram_data_T_224_en;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  T_221;
  wire  T_222;
  wire  do_enq;
  wire  T_223;
  wire  do_deq;
  wire  T_249;
  wire  GEN_17;
  wire  T_251;
  wire [1:0] T_277;
  wire  ptr_diff;
  wire [1:0] T_279;
  assign io_enq_ready = T_221;
  assign io_deq_valid = T_251;
  assign io_deq_bits_addr_block = ram_addr_block_T_254_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_254_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_254_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_254_data;
  assign io_deq_bits_a_type = ram_a_type_T_254_data;
  assign io_deq_bits_union = ram_union_T_254_data;
  assign io_deq_bits_data = ram_data_T_254_data;
  assign io_count = T_279[0];
  assign ram_addr_block_T_254_addr = 1'h0;
  assign ram_addr_block_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_block_T_254_data = ram_addr_block[ram_addr_block_T_254_addr];
  `else
  assign ram_addr_block_T_254_data = ram_addr_block_T_254_addr >= 1'h1 ? $random : ram_addr_block[ram_addr_block_T_254_addr];
  `endif
  assign ram_addr_block_T_224_data = io_enq_bits_addr_block;
  assign ram_addr_block_T_224_addr = 1'h0;
  assign ram_addr_block_T_224_mask = do_enq;
  assign ram_addr_block_T_224_en = do_enq;
  assign ram_client_xact_id_T_254_addr = 1'h0;
  assign ram_client_xact_id_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_client_xact_id_T_254_data = ram_client_xact_id[ram_client_xact_id_T_254_addr];
  `else
  assign ram_client_xact_id_T_254_data = ram_client_xact_id_T_254_addr >= 1'h1 ? $random : ram_client_xact_id[ram_client_xact_id_T_254_addr];
  `endif
  assign ram_client_xact_id_T_224_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_224_addr = 1'h0;
  assign ram_client_xact_id_T_224_mask = do_enq;
  assign ram_client_xact_id_T_224_en = do_enq;
  assign ram_addr_beat_T_254_addr = 1'h0;
  assign ram_addr_beat_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_beat_T_254_data = ram_addr_beat[ram_addr_beat_T_254_addr];
  `else
  assign ram_addr_beat_T_254_data = ram_addr_beat_T_254_addr >= 1'h1 ? $random : ram_addr_beat[ram_addr_beat_T_254_addr];
  `endif
  assign ram_addr_beat_T_224_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_224_addr = 1'h0;
  assign ram_addr_beat_T_224_mask = do_enq;
  assign ram_addr_beat_T_224_en = do_enq;
  assign ram_is_builtin_type_T_254_addr = 1'h0;
  assign ram_is_builtin_type_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_is_builtin_type_T_254_data = ram_is_builtin_type[ram_is_builtin_type_T_254_addr];
  `else
  assign ram_is_builtin_type_T_254_data = ram_is_builtin_type_T_254_addr >= 1'h1 ? $random : ram_is_builtin_type[ram_is_builtin_type_T_254_addr];
  `endif
  assign ram_is_builtin_type_T_224_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_224_addr = 1'h0;
  assign ram_is_builtin_type_T_224_mask = do_enq;
  assign ram_is_builtin_type_T_224_en = do_enq;
  assign ram_a_type_T_254_addr = 1'h0;
  assign ram_a_type_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_a_type_T_254_data = ram_a_type[ram_a_type_T_254_addr];
  `else
  assign ram_a_type_T_254_data = ram_a_type_T_254_addr >= 1'h1 ? $random : ram_a_type[ram_a_type_T_254_addr];
  `endif
  assign ram_a_type_T_224_data = io_enq_bits_a_type;
  assign ram_a_type_T_224_addr = 1'h0;
  assign ram_a_type_T_224_mask = do_enq;
  assign ram_a_type_T_224_en = do_enq;
  assign ram_union_T_254_addr = 1'h0;
  assign ram_union_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_union_T_254_data = ram_union[ram_union_T_254_addr];
  `else
  assign ram_union_T_254_data = ram_union_T_254_addr >= 1'h1 ? $random : ram_union[ram_union_T_254_addr];
  `endif
  assign ram_union_T_224_data = io_enq_bits_union;
  assign ram_union_T_224_addr = 1'h0;
  assign ram_union_T_224_mask = do_enq;
  assign ram_union_T_224_en = do_enq;
  assign ram_data_T_254_addr = 1'h0;
  assign ram_data_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_data_T_254_data = ram_data[ram_data_T_254_addr];
  `else
  assign ram_data_T_254_data = ram_data_T_254_addr >= 1'h1 ? $random : ram_data[ram_data_T_254_addr];
  `endif
  assign ram_data_T_224_data = io_enq_bits_data;
  assign ram_data_T_224_addr = 1'h0;
  assign ram_data_T_224_mask = do_enq;
  assign ram_data_T_224_en = do_enq;
  assign T_221 = maybe_full == 1'h0;
  assign T_222 = io_enq_ready & io_enq_valid;
  assign do_enq = T_222;
  assign T_223 = io_deq_ready & io_deq_valid;
  assign do_deq = T_223;
  assign T_249 = do_enq != do_deq;
  assign GEN_17 = T_249 ? do_enq : maybe_full;
  assign T_251 = T_221 == 1'h0;
  assign T_277 = 1'h0 - 1'h0;
  assign ptr_diff = T_277[0:0];
  assign T_279 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_block[initvar] = GEN_0[25:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[1:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_2[2:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_union[initvar] = GEN_5[11:0];
  GEN_6 = {2{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_6[63:0];
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_block_T_224_en & ram_addr_block_T_224_mask) begin
      ram_addr_block[ram_addr_block_T_224_addr] <= ram_addr_block_T_224_data;
    end
    if(ram_client_xact_id_T_224_en & ram_client_xact_id_T_224_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_224_addr] <= ram_client_xact_id_T_224_data;
    end
    if(ram_addr_beat_T_224_en & ram_addr_beat_T_224_mask) begin
      ram_addr_beat[ram_addr_beat_T_224_addr] <= ram_addr_beat_T_224_data;
    end
    if(ram_is_builtin_type_T_224_en & ram_is_builtin_type_T_224_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_224_addr] <= ram_is_builtin_type_T_224_data;
    end
    if(ram_a_type_T_224_en & ram_a_type_T_224_mask) begin
      ram_a_type[ram_a_type_T_224_addr] <= ram_a_type_T_224_data;
    end
    if(ram_union_T_224_en & ram_union_T_224_mask) begin
      ram_union[ram_union_T_224_addr] <= ram_union_T_224_data;
    end
    if(ram_data_T_224_en & ram_data_T_224_mask) begin
      ram_data[ram_data_T_224_addr] <= ram_data_T_224_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_249) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module PLIC(
  input   clk,
  input   reset,
  input   io_devices_0_valid,
  output  io_devices_0_ready,
  output  io_devices_0_complete,
  input   io_devices_1_valid,
  output  io_devices_1_ready,
  output  io_devices_1_complete,
  output  io_harts_0,
  output  io_harts_1,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data
);
  wire  T_477_0;
  wire  T_477_1;
  wire  T_477_2;
  wire  priority_0;
  wire  priority_1;
  wire  priority_2;
  wire  T_489_0;
  wire  T_489_1;
  wire  threshold_0;
  wire  threshold_1;
  wire  T_502_0;
  wire  T_502_1;
  wire  T_502_2;
  reg  pending_0;
  reg [31:0] GEN_15;
  reg  pending_1;
  reg [31:0] GEN_18;
  reg  pending_2;
  reg [31:0] GEN_19;
  reg  enables_0_0;
  reg [31:0] GEN_29;
  reg  enables_0_1;
  reg [31:0] GEN_32;
  reg  enables_0_2;
  reg [31:0] GEN_33;
  reg  enables_1_0;
  reg [31:0] GEN_36;
  reg  enables_1_1;
  reg [31:0] GEN_37;
  reg  enables_1_2;
  reg [31:0] GEN_38;
  wire  T_545;
  wire  GEN_11;
  wire  T_549;
  wire  GEN_12;
  wire [1:0] maxDevs_0;
  wire [1:0] maxDevs_1;
  wire  T_559;
  wire [1:0] T_560;
  wire  T_561;
  wire [1:0] T_562;
  wire  T_567;
  wire [1:0] T_568;
  wire [1:0] T_570;
  wire  T_571;
  wire  T_572;
  wire  T_574;
  wire [1:0] T_575;
  wire [1:0] GEN_101;
  wire [2:0] T_577;
  wire [1:0] T_578;
  wire [1:0] T_579;
  reg [1:0] T_580;
  reg [31:0] GEN_41;
  reg [1:0] T_581;
  reg [31:0] GEN_43;
  wire [1:0] T_583;
  wire  T_584;
  wire  T_585;
  wire [1:0] T_586;
  wire  T_587;
  wire [1:0] T_588;
  wire  T_593;
  wire [1:0] T_594;
  wire  T_598;
  wire  T_600;
  wire [1:0] T_601;
  wire [1:0] T_605;
  reg [1:0] T_606;
  reg [31:0] GEN_44;
  reg [1:0] T_607;
  reg [31:0] GEN_47;
  wire [1:0] T_609;
  wire  T_610;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_634;
  wire  T_636;
  wire  T_637;
  wire  read;
  wire  T_640;
  wire  T_641;
  wire  write;
  wire  T_644;
  wire  T_645;
  wire  T_646;
  wire  T_647;
  wire  T_649;
  wire [2:0] T_650;
  wire [28:0] T_651;
  wire [31:0] T_652;
  wire [25:0] addr;
  wire [25:0] GEN_103;
  wire [26:0] T_654;
  wire [25:0] T_655;
  wire  claimant;
  wire  hart;
  wire [1:0] GEN_0;
  wire [1:0] GEN_13;
  wire [2:0] T_657;
  wire [1:0] myMaxDev;
  wire [63:0] rdata;
  wire  T_663;
  wire  T_664;
  wire [7:0] GEN_105;
  wire [8:0] T_668;
  wire [7:0] T_669;
  wire [7:0] T_675_0;
  wire  T_678;
  wire  T_679;
  wire  T_683;
  wire [7:0] T_684;
  wire [7:0] T_686;
  wire [7:0] T_687;
  wire  T_688;
  wire  T_689;
  wire  T_690;
  wire  T_691;
  wire  T_692;
  wire  T_693;
  wire  T_694;
  wire  T_695;
  wire [7:0] GEN_106;
  wire [8:0] T_697;
  wire [7:0] T_698;
  wire [7:0] GEN_107;
  wire [8:0] T_700;
  wire [7:0] T_701;
  wire [7:0] GEN_108;
  wire [8:0] T_703;
  wire [7:0] T_704;
  wire [7:0] GEN_109;
  wire [8:0] T_706;
  wire [7:0] T_707;
  wire [7:0] GEN_110;
  wire [8:0] T_709;
  wire [7:0] T_710;
  wire [7:0] GEN_111;
  wire [8:0] T_712;
  wire [7:0] T_713;
  wire [7:0] GEN_112;
  wire [8:0] T_715;
  wire [7:0] T_716;
  wire [7:0] GEN_113;
  wire [8:0] T_718;
  wire [7:0] T_719;
  wire [7:0] T_725_0;
  wire [7:0] T_725_1;
  wire [7:0] T_725_2;
  wire [7:0] T_725_3;
  wire [7:0] T_725_4;
  wire [7:0] T_725_5;
  wire [7:0] T_725_6;
  wire [7:0] T_725_7;
  wire [15:0] T_727;
  wire [15:0] T_728;
  wire [31:0] T_729;
  wire [15:0] T_730;
  wire [15:0] T_731;
  wire [31:0] T_732;
  wire [63:0] T_733;
  wire [63:0] T_734;
  wire [7:0] T_748_0;
  wire [7:0] T_760;
  wire  T_761;
  wire  T_762;
  wire  T_763;
  wire  T_764;
  wire  T_765;
  wire  T_766;
  wire  T_767;
  wire  T_768;
  wire [7:0] GEN_115;
  wire [8:0] T_770;
  wire [7:0] T_771;
  wire [7:0] GEN_116;
  wire [8:0] T_773;
  wire [7:0] T_774;
  wire [7:0] GEN_117;
  wire [8:0] T_776;
  wire [7:0] T_777;
  wire [7:0] GEN_118;
  wire [8:0] T_779;
  wire [7:0] T_780;
  wire [7:0] GEN_119;
  wire [8:0] T_782;
  wire [7:0] T_783;
  wire [7:0] GEN_120;
  wire [8:0] T_785;
  wire [7:0] T_786;
  wire [7:0] GEN_121;
  wire [8:0] T_788;
  wire [7:0] T_789;
  wire [7:0] GEN_122;
  wire [8:0] T_791;
  wire [7:0] T_792;
  wire [7:0] T_798_0;
  wire [7:0] T_798_1;
  wire [7:0] T_798_2;
  wire [7:0] T_798_3;
  wire [7:0] T_798_4;
  wire [7:0] T_798_5;
  wire [7:0] T_798_6;
  wire [7:0] T_798_7;
  wire [15:0] T_800;
  wire [15:0] T_801;
  wire [31:0] T_802;
  wire [15:0] T_803;
  wire [15:0] T_804;
  wire [31:0] T_805;
  wire [63:0] T_806;
  wire [63:0] T_807;
  wire [63:0] T_808;
  wire [63:0] masked_wdata;
  wire  T_810;
  wire [32:0] T_813;
  wire  GEN_1;
  wire  GEN_14;
  wire [33:0] T_814;
  wire [6:0] GEN_124;
  wire [7:0] T_816;
  wire [33:0] T_817;
  wire  T_818;
  wire  T_819;
  wire  GEN_2;
  wire [1:0] GEN_126;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_20;
  wire  GEN_21;
  wire [7:0] T_834_0;
  wire [7:0] T_846;
  wire  T_847;
  wire [31:0] T_848;
  wire [1:0] T_849;
  wire  GEN_3;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_22;
  wire  GEN_132;
  wire  GEN_23;
  wire  GEN_134;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire [2:0] T_851;
  wire [1:0] T_852;
  wire  GEN_4;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_39;
  wire  GEN_40;
  wire [63:0] GEN_42;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_50;
  wire  GEN_51;
  wire [25:0] GEN_141;
  wire  T_860;
  wire  T_862;
  wire  T_863;
  wire [26:0] T_865;
  wire [25:0] T_866;
  wire  T_867;
  wire  GEN_5;
  wire  GEN_52;
  wire  GEN_6;
  wire  GEN_53;
  wire [1:0] T_871;
  wire  GEN_7;
  wire  GEN_54;
  wire [2:0] T_872;
  wire  T_876;
  wire  GEN_8;
  wire  T_880;
  wire  GEN_9;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_63;
  wire  GEN_64;
  wire  T_884;
  wire  GEN_10;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_68;
  wire  GEN_69;
  wire [63:0] GEN_73;
  wire  GEN_83;
  wire [63:0] GEN_87;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_95;
  wire  GEN_96;
  wire [25:0] GEN_143;
  wire  T_886;
  wire  T_890;
  wire  T_891;
  wire  T_892;
  wire [1:0] T_894;
  wire [2:0] T_895;
  wire [2:0] T_898;
  wire [63:0] GEN_97;
  wire  T_905;
  wire  T_906;
  wire  T_907;
  wire  T_909;
  wire [31:0] T_911;
  wire [31:0] T_913;
  wire [63:0] T_914;
  wire [63:0] GEN_98;
  wire [31:0] T_918;
  wire [63:0] GEN_99;
  wire [63:0] GEN_100;
  wire  T_939;
  wire [2:0] T_940;
  wire  T_941;
  wire [2:0] T_942;
  wire  T_943;
  wire [2:0] T_944;
  wire  T_945;
  wire [2:0] T_946;
  wire  T_947;
  wire [2:0] T_948;
  wire  T_949;
  wire [2:0] T_950;
  wire  T_951;
  wire [2:0] T_952;
  wire [2:0] T_977_addr_beat;
  wire [1:0] T_977_client_xact_id;
  wire  T_977_manager_xact_id;
  wire  T_977_is_builtin_type;
  wire [3:0] T_977_g_type;
  wire [63:0] T_977_data;
  Queue_20 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_devices_0_ready = T_545;
  assign io_devices_0_complete = GEN_50;
  assign io_devices_1_ready = T_549;
  assign io_devices_1_complete = GEN_51;
  assign io_harts_0 = T_584;
  assign io_harts_1 = T_610;
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_977_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_977_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_977_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_977_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_977_g_type;
  assign io_tl_grant_bits_data = T_977_data;
  assign T_477_0 = 1'h1;
  assign T_477_1 = 1'h1;
  assign T_477_2 = 1'h1;
  assign priority_0 = 1'h0;
  assign priority_1 = T_477_1;
  assign priority_2 = T_477_2;
  assign T_489_0 = 1'h0;
  assign T_489_1 = 1'h0;
  assign threshold_0 = T_489_0;
  assign threshold_1 = T_489_1;
  assign T_502_0 = 1'h0;
  assign T_502_1 = 1'h0;
  assign T_502_2 = 1'h0;
  assign T_545 = pending_1 == 1'h0;
  assign GEN_11 = io_devices_0_valid ? 1'h1 : pending_1;
  assign T_549 = pending_2 == 1'h0;
  assign GEN_12 = io_devices_1_valid ? 1'h1 : pending_2;
  assign maxDevs_0 = T_580;
  assign maxDevs_1 = T_606;
  assign T_559 = pending_1 & enables_0_1;
  assign T_560 = {T_559,priority_1};
  assign T_561 = pending_2 & enables_0_2;
  assign T_562 = {T_561,priority_2};
  assign T_567 = 2'h2 >= T_560;
  assign T_568 = T_567 ? 2'h2 : T_560;
  assign T_570 = 1'h1 + 1'h0;
  assign T_571 = T_570[0:0];
  assign T_572 = T_567 ? 1'h0 : T_571;
  assign T_574 = T_568 >= T_562;
  assign T_575 = T_574 ? T_568 : T_562;
  assign GEN_101 = {{1'd0}, 1'h0};
  assign T_577 = 2'h2 + GEN_101;
  assign T_578 = T_577[1:0];
  assign T_579 = T_574 ? {{1'd0}, T_572} : T_578;
  assign T_583 = {1'h1,threshold_0};
  assign T_584 = T_581 > T_583;
  assign T_585 = pending_1 & enables_1_1;
  assign T_586 = {T_585,priority_1};
  assign T_587 = pending_2 & enables_1_2;
  assign T_588 = {T_587,priority_2};
  assign T_593 = 2'h2 >= T_586;
  assign T_594 = T_593 ? 2'h2 : T_586;
  assign T_598 = T_593 ? 1'h0 : T_571;
  assign T_600 = T_594 >= T_588;
  assign T_601 = T_600 ? T_594 : T_588;
  assign T_605 = T_600 ? {{1'd0}, T_598} : T_578;
  assign T_609 = {1'h1,threshold_1};
  assign T_610 = T_607 > T_609;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_634 = acq_io_deq_ready & acq_io_deq_valid;
  assign T_636 = acq_io_deq_bits_a_type == 3'h0;
  assign T_637 = acq_io_deq_bits_is_builtin_type & T_636;
  assign read = T_634 & T_637;
  assign T_640 = acq_io_deq_bits_a_type == 3'h2;
  assign T_641 = acq_io_deq_bits_is_builtin_type & T_640;
  assign write = T_634 & T_641;
  assign T_644 = T_634 == 1'h0;
  assign T_645 = T_644 | read;
  assign T_646 = T_645 | write;
  assign T_647 = T_646 | reset;
  assign T_649 = T_647 == 1'h0;
  assign T_650 = acq_io_deq_bits_union[11:9];
  assign T_651 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_652 = {T_651,T_650};
  assign addr = T_652[25:0];
  assign GEN_103 = {{4'd0}, 22'h200000};
  assign T_654 = addr - GEN_103;
  assign T_655 = T_654[25:0];
  assign claimant = T_655[12];
  assign hart = GEN_83;
  assign GEN_0 = GEN_13;
  assign GEN_13 = claimant ? maxDevs_1 : maxDevs_0;
  assign T_657 = GEN_0 + GEN_101;
  assign myMaxDev = T_657[1:0];
  assign rdata = GEN_100;
  assign T_663 = acq_io_deq_bits_a_type == 3'h4;
  assign T_664 = acq_io_deq_bits_is_builtin_type & T_663;
  assign GEN_105 = {{7'd0}, 1'h1};
  assign T_668 = 8'h0 - GEN_105;
  assign T_669 = T_668[7:0];
  assign T_675_0 = T_669;
  assign T_678 = acq_io_deq_bits_a_type == 3'h3;
  assign T_679 = acq_io_deq_bits_is_builtin_type & T_678;
  assign T_683 = T_679 | T_641;
  assign T_684 = acq_io_deq_bits_union[8:1];
  assign T_686 = T_683 ? T_684 : {{7'd0}, 1'h0};
  assign T_687 = T_664 ? T_675_0 : T_686;
  assign T_688 = T_687[0];
  assign T_689 = T_687[1];
  assign T_690 = T_687[2];
  assign T_691 = T_687[3];
  assign T_692 = T_687[4];
  assign T_693 = T_687[5];
  assign T_694 = T_687[6];
  assign T_695 = T_687[7];
  assign GEN_106 = {{7'd0}, T_688};
  assign T_697 = 8'h0 - GEN_106;
  assign T_698 = T_697[7:0];
  assign GEN_107 = {{7'd0}, T_689};
  assign T_700 = 8'h0 - GEN_107;
  assign T_701 = T_700[7:0];
  assign GEN_108 = {{7'd0}, T_690};
  assign T_703 = 8'h0 - GEN_108;
  assign T_704 = T_703[7:0];
  assign GEN_109 = {{7'd0}, T_691};
  assign T_706 = 8'h0 - GEN_109;
  assign T_707 = T_706[7:0];
  assign GEN_110 = {{7'd0}, T_692};
  assign T_709 = 8'h0 - GEN_110;
  assign T_710 = T_709[7:0];
  assign GEN_111 = {{7'd0}, T_693};
  assign T_712 = 8'h0 - GEN_111;
  assign T_713 = T_712[7:0];
  assign GEN_112 = {{7'd0}, T_694};
  assign T_715 = 8'h0 - GEN_112;
  assign T_716 = T_715[7:0];
  assign GEN_113 = {{7'd0}, T_695};
  assign T_718 = 8'h0 - GEN_113;
  assign T_719 = T_718[7:0];
  assign T_725_0 = T_698;
  assign T_725_1 = T_701;
  assign T_725_2 = T_704;
  assign T_725_3 = T_707;
  assign T_725_4 = T_710;
  assign T_725_5 = T_713;
  assign T_725_6 = T_716;
  assign T_725_7 = T_719;
  assign T_727 = {T_725_1,T_725_0};
  assign T_728 = {T_725_3,T_725_2};
  assign T_729 = {T_728,T_727};
  assign T_730 = {T_725_5,T_725_4};
  assign T_731 = {T_725_7,T_725_6};
  assign T_732 = {T_731,T_730};
  assign T_733 = {T_732,T_729};
  assign T_734 = acq_io_deq_bits_data & T_733;
  assign T_748_0 = T_669;
  assign T_760 = T_664 ? T_748_0 : T_686;
  assign T_761 = T_760[0];
  assign T_762 = T_760[1];
  assign T_763 = T_760[2];
  assign T_764 = T_760[3];
  assign T_765 = T_760[4];
  assign T_766 = T_760[5];
  assign T_767 = T_760[6];
  assign T_768 = T_760[7];
  assign GEN_115 = {{7'd0}, T_761};
  assign T_770 = 8'h0 - GEN_115;
  assign T_771 = T_770[7:0];
  assign GEN_116 = {{7'd0}, T_762};
  assign T_773 = 8'h0 - GEN_116;
  assign T_774 = T_773[7:0];
  assign GEN_117 = {{7'd0}, T_763};
  assign T_776 = 8'h0 - GEN_117;
  assign T_777 = T_776[7:0];
  assign GEN_118 = {{7'd0}, T_764};
  assign T_779 = 8'h0 - GEN_118;
  assign T_780 = T_779[7:0];
  assign GEN_119 = {{7'd0}, T_765};
  assign T_782 = 8'h0 - GEN_119;
  assign T_783 = T_782[7:0];
  assign GEN_120 = {{7'd0}, T_766};
  assign T_785 = 8'h0 - GEN_120;
  assign T_786 = T_785[7:0];
  assign GEN_121 = {{7'd0}, T_767};
  assign T_788 = 8'h0 - GEN_121;
  assign T_789 = T_788[7:0];
  assign GEN_122 = {{7'd0}, T_768};
  assign T_791 = 8'h0 - GEN_122;
  assign T_792 = T_791[7:0];
  assign T_798_0 = T_771;
  assign T_798_1 = T_774;
  assign T_798_2 = T_777;
  assign T_798_3 = T_780;
  assign T_798_4 = T_783;
  assign T_798_5 = T_786;
  assign T_798_6 = T_789;
  assign T_798_7 = T_792;
  assign T_800 = {T_798_1,T_798_0};
  assign T_801 = {T_798_3,T_798_2};
  assign T_802 = {T_801,T_800};
  assign T_803 = {T_798_5,T_798_4};
  assign T_804 = {T_798_7,T_798_6};
  assign T_805 = {T_804,T_803};
  assign T_806 = {T_805,T_802};
  assign T_807 = ~ T_806;
  assign T_808 = rdata & T_807;
  assign masked_wdata = T_734 | T_808;
  assign T_810 = addr >= GEN_103;
  assign T_813 = {myMaxDev,31'h0};
  assign GEN_1 = GEN_14;
  assign GEN_14 = claimant ? threshold_1 : threshold_0;
  assign T_814 = {T_813,GEN_1};
  assign GEN_124 = {{6'd0}, 1'h0};
  assign T_816 = GEN_124 * 7'h40;
  assign T_817 = T_814 >> T_816;
  assign T_818 = addr[2];
  assign T_819 = read & T_818;
  assign GEN_2 = 1'h0;
  assign GEN_126 = {{1'd0}, 1'h1};
  assign GEN_16 = GEN_126 == myMaxDev ? GEN_2 : GEN_11;
  assign GEN_17 = 2'h2 == myMaxDev ? GEN_2 : GEN_12;
  assign GEN_20 = T_819 ? GEN_16 : GEN_11;
  assign GEN_21 = T_819 ? GEN_17 : GEN_12;
  assign T_834_0 = T_669;
  assign T_846 = T_664 ? T_834_0 : T_686;
  assign T_847 = T_846[4];
  assign T_848 = acq_io_deq_bits_data[63:32];
  assign T_849 = T_848[1:0];
  assign GEN_3 = GEN_26;
  assign GEN_129 = 1'h0 == hart;
  assign GEN_130 = GEN_126 == T_849;
  assign GEN_22 = GEN_129 & GEN_130 ? enables_0_1 : enables_0_0;
  assign GEN_132 = 2'h2 == T_849;
  assign GEN_23 = GEN_129 & GEN_132 ? enables_0_2 : GEN_22;
  assign GEN_134 = GEN_101 == T_849;
  assign GEN_24 = hart & GEN_134 ? enables_1_0 : GEN_23;
  assign GEN_25 = hart & GEN_130 ? enables_1_1 : GEN_24;
  assign GEN_26 = hart & GEN_132 ? enables_1_2 : GEN_25;
  assign T_851 = T_849 - GEN_126;
  assign T_852 = T_851[1:0];
  assign GEN_4 = 1'h1;
  assign GEN_27 = GEN_101 == T_852 ? GEN_4 : 1'h0;
  assign GEN_28 = GEN_126 == T_852 ? GEN_4 : 1'h0;
  assign GEN_30 = GEN_3 ? GEN_27 : 1'h0;
  assign GEN_31 = GEN_3 ? GEN_28 : 1'h0;
  assign GEN_34 = T_847 ? GEN_30 : 1'h0;
  assign GEN_35 = T_847 ? GEN_31 : 1'h0;
  assign GEN_39 = write ? GEN_34 : 1'h0;
  assign GEN_40 = write ? GEN_35 : 1'h0;
  assign GEN_42 = T_810 ? {{30'd0}, T_817} : 64'h0;
  assign GEN_45 = T_810 ? GEN_20 : GEN_11;
  assign GEN_46 = T_810 ? GEN_21 : GEN_12;
  assign GEN_50 = T_810 ? GEN_39 : 1'h0;
  assign GEN_51 = T_810 ? GEN_40 : 1'h0;
  assign GEN_141 = {{12'd0}, 14'h2000};
  assign T_860 = addr >= GEN_141;
  assign T_862 = T_810 == 1'h0;
  assign T_863 = T_862 & T_860;
  assign T_865 = addr - GEN_141;
  assign T_866 = T_865[25:0];
  assign T_867 = T_866[7];
  assign GEN_5 = GEN_52;
  assign GEN_52 = hart ? enables_1_2 : enables_0_2;
  assign GEN_6 = GEN_53;
  assign GEN_53 = hart ? enables_1_1 : enables_0_1;
  assign T_871 = {GEN_5,GEN_6};
  assign GEN_7 = GEN_54;
  assign GEN_54 = hart ? enables_1_0 : enables_0_0;
  assign T_872 = {T_871,GEN_7};
  assign T_876 = masked_wdata[0];
  assign GEN_8 = T_876;
  assign T_880 = masked_wdata[1];
  assign GEN_9 = T_880;
  assign GEN_60 = 1'h0 == T_867 ? GEN_9 : enables_0_1;
  assign GEN_61 = T_867 ? GEN_9 : enables_1_1;
  assign GEN_63 = write ? GEN_60 : enables_0_1;
  assign GEN_64 = write ? GEN_61 : enables_1_1;
  assign T_884 = masked_wdata[2];
  assign GEN_10 = T_884;
  assign GEN_65 = 1'h0 == T_867 ? GEN_10 : enables_0_2;
  assign GEN_66 = T_867 ? GEN_10 : enables_1_2;
  assign GEN_68 = write ? GEN_65 : enables_0_2;
  assign GEN_69 = write ? GEN_66 : enables_1_2;
  assign GEN_73 = 1'h1 ? {{61'd0}, T_872} : GEN_42;
  assign GEN_83 = T_863 ? T_867 : claimant;
  assign GEN_87 = T_863 ? GEN_73 : GEN_42;
  assign GEN_92 = T_863 ? GEN_63 : enables_0_1;
  assign GEN_93 = T_863 ? GEN_64 : enables_1_1;
  assign GEN_95 = T_863 ? GEN_68 : enables_0_2;
  assign GEN_96 = T_863 ? GEN_69 : enables_1_2;
  assign GEN_143 = {{13'd0}, 13'h1000};
  assign T_886 = addr >= GEN_143;
  assign T_890 = T_860 == 1'h0;
  assign T_891 = T_862 & T_890;
  assign T_892 = T_891 & T_886;
  assign T_894 = {pending_2,pending_1};
  assign T_895 = {T_894,pending_0};
  assign T_898 = T_895 >> T_816;
  assign GEN_97 = T_892 ? {{61'd0}, T_898} : GEN_87;
  assign T_905 = T_886 == 1'h0;
  assign T_906 = T_891 & T_905;
  assign T_907 = addr[3];
  assign T_909 = T_907 == 1'h0;
  assign T_911 = {31'h0,priority_0};
  assign T_913 = {31'h0,priority_1};
  assign T_914 = {T_913,T_911};
  assign GEN_98 = T_909 ? T_914 : GEN_97;
  assign T_918 = {31'h0,priority_2};
  assign GEN_99 = T_907 ? {{32'd0}, T_918} : GEN_98;
  assign GEN_100 = T_906 ? GEN_99 : GEN_97;
  assign T_939 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_940 = T_939 ? 3'h1 : 3'h3;
  assign T_941 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_942 = T_941 ? 3'h1 : T_940;
  assign T_943 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_944 = T_943 ? 3'h4 : T_942;
  assign T_945 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_946 = T_945 ? 3'h3 : T_944;
  assign T_947 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_948 = T_947 ? 3'h3 : T_946;
  assign T_949 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_950 = T_949 ? 3'h5 : T_948;
  assign T_951 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_952 = T_951 ? 3'h4 : T_950;
  assign T_977_addr_beat = {{2'd0}, 1'h0};
  assign T_977_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_977_manager_xact_id = 1'h0;
  assign T_977_is_builtin_type = 1'h1;
  assign T_977_g_type = {{1'd0}, T_952};
  assign T_977_data = rdata;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  pending_0 = GEN_15[0:0];
  GEN_18 = {1{$random}};
  pending_1 = GEN_18[0:0];
  GEN_19 = {1{$random}};
  pending_2 = GEN_19[0:0];
  GEN_29 = {1{$random}};
  enables_0_0 = GEN_29[0:0];
  GEN_32 = {1{$random}};
  enables_0_1 = GEN_32[0:0];
  GEN_33 = {1{$random}};
  enables_0_2 = GEN_33[0:0];
  GEN_36 = {1{$random}};
  enables_1_0 = GEN_36[0:0];
  GEN_37 = {1{$random}};
  enables_1_1 = GEN_37[0:0];
  GEN_38 = {1{$random}};
  enables_1_2 = GEN_38[0:0];
  GEN_41 = {1{$random}};
  T_580 = GEN_41[1:0];
  GEN_43 = {1{$random}};
  T_581 = GEN_43[1:0];
  GEN_44 = {1{$random}};
  T_606 = GEN_44[1:0];
  GEN_47 = {1{$random}};
  T_607 = GEN_47[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      pending_0 <= T_502_0;
    end else begin
      pending_0 <= 1'h0;
    end
    if(reset) begin
      pending_1 <= T_502_1;
    end else begin
      if(T_810) begin
        if(T_819) begin
          if(GEN_126 == myMaxDev) begin
            pending_1 <= GEN_2;
          end else begin
            if(io_devices_0_valid) begin
              pending_1 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_0_valid) begin
            pending_1 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_0_valid) begin
          pending_1 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_2 <= T_502_2;
    end else begin
      if(T_810) begin
        if(T_819) begin
          if(2'h2 == myMaxDev) begin
            pending_2 <= GEN_2;
          end else begin
            if(io_devices_1_valid) begin
              pending_2 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_1_valid) begin
            pending_2 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_1_valid) begin
          pending_2 <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      enables_0_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(T_863) begin
        if(write) begin
          if(1'h0 == T_867) begin
            enables_0_1 <= GEN_9;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_863) begin
        if(write) begin
          if(1'h0 == T_867) begin
            enables_0_2 <= GEN_10;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      enables_1_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(T_863) begin
        if(write) begin
          if(T_867) begin
            enables_1_1 <= GEN_9;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_863) begin
        if(write) begin
          if(T_867) begin
            enables_1_2 <= GEN_10;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_574) begin
        T_580 <= {{1'd0}, T_572};
      end else begin
        T_580 <= T_578;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_574) begin
        if(T_567) begin
          T_581 <= 2'h2;
        end else begin
          T_581 <= T_560;
        end
      end else begin
        T_581 <= T_562;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_600) begin
        T_606 <= {{1'd0}, T_598};
      end else begin
        T_606 <= T_578;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_600) begin
        if(T_593) begin
          T_607 <= 2'h2;
        end else begin
          T_607 <= T_586;
        end
      end else begin
        T_607 <= T_588;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_649) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported PLIC operation\n    at Plic.scala:108 assert(!acq.fire() || read || write, \"unsupported PLIC operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_649) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_649) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module LevelGateway(
  input   clk,
  input   reset,
  input   io_interrupt,
  output  io_plic_valid,
  input   io_plic_ready,
  input   io_plic_complete
);
  reg  inFlight;
  reg [31:0] GEN_2;
  wire  T_6;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_10;
  wire  T_11;
  assign io_plic_valid = T_11;
  assign T_6 = io_interrupt & io_plic_ready;
  assign GEN_0 = T_6 ? 1'h1 : inFlight;
  assign GEN_1 = io_plic_complete ? 1'h0 : GEN_0;
  assign T_10 = inFlight == 1'h0;
  assign T_11 = io_interrupt & T_10;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_2 = {1{$random}};
  inFlight = GEN_2[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      inFlight <= 1'h0;
    end else begin
      if(io_plic_complete) begin
        inFlight <= 1'h0;
      end else begin
        if(T_6) begin
          inFlight <= 1'h1;
        end
      end
    end
  end
endmodule
module DebugModule(
  input   clk,
  input   reset,
  output  io_db_req_ready,
  input   io_db_req_valid,
  input  [4:0] io_db_req_bits_addr,
  input  [1:0] io_db_req_bits_op,
  input  [33:0] io_db_req_bits_data,
  input   io_db_resp_ready,
  output  io_db_resp_valid,
  output [1:0] io_db_resp_bits_resp,
  output [33:0] io_db_resp_bits_data,
  output  io_debugInterrupts_0,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_ndreset,
  output  io_fullreset
);
  wire  CONTROLReset_interrupt;
  wire  CONTROLReset_haltnot;
  wire [9:0] CONTROLReset_reserved0;
  wire [2:0] CONTROLReset_buserror;
  wire [2:0] CONTROLReset_serial;
  wire  CONTROLReset_autoincrement;
  wire [2:0] CONTROLReset_access;
  wire [9:0] CONTROLReset_hartid;
  wire  CONTROLReset_ndreset;
  wire  CONTROLReset_fullreset;
  wire  CONTROLWrEn;
  reg  CONTROLReg_interrupt;
  reg [31:0] GEN_26;
  reg  CONTROLReg_haltnot;
  reg [31:0] GEN_27;
  reg [9:0] CONTROLReg_reserved0;
  reg [31:0] GEN_28;
  reg [2:0] CONTROLReg_buserror;
  reg [31:0] GEN_29;
  reg [2:0] CONTROLReg_serial;
  reg [31:0] GEN_30;
  reg  CONTROLReg_autoincrement;
  reg [31:0] GEN_52;
  reg [2:0] CONTROLReg_access;
  reg [31:0] GEN_85;
  reg [9:0] CONTROLReg_hartid;
  reg [31:0] GEN_86;
  reg  CONTROLReg_ndreset;
  reg [31:0] GEN_88;
  reg  CONTROLReg_fullreset;
  reg [31:0] GEN_89;
  wire  CONTROLWrData_interrupt;
  wire  CONTROLWrData_haltnot;
  wire [9:0] CONTROLWrData_reserved0;
  wire [2:0] CONTROLWrData_buserror;
  wire [2:0] CONTROLWrData_serial;
  wire  CONTROLWrData_autoincrement;
  wire [2:0] CONTROLWrData_access;
  wire [9:0] CONTROLWrData_hartid;
  wire  CONTROLWrData_ndreset;
  wire  CONTROLWrData_fullreset;
  wire  CONTROLRdData_interrupt;
  wire  CONTROLRdData_haltnot;
  wire [9:0] CONTROLRdData_reserved0;
  wire [2:0] CONTROLRdData_buserror;
  wire [2:0] CONTROLRdData_serial;
  wire  CONTROLRdData_autoincrement;
  wire [2:0] CONTROLRdData_access;
  wire [9:0] CONTROLRdData_hartid;
  wire  CONTROLRdData_ndreset;
  wire  CONTROLRdData_fullreset;
  reg  ndresetCtrReg;
  reg [31:0] GEN_90;
  wire [1:0] DMINFORdData_reserved0;
  wire [6:0] DMINFORdData_abussize;
  wire [3:0] DMINFORdData_serialcount;
  wire  DMINFORdData_access128;
  wire  DMINFORdData_access64;
  wire  DMINFORdData_access32;
  wire  DMINFORdData_access16;
  wire  DMINFORdData_accesss8;
  wire [5:0] DMINFORdData_dramsize;
  wire  DMINFORdData_haltsum;
  wire [2:0] DMINFORdData_reserved1;
  wire  DMINFORdData_authenticated;
  wire  DMINFORdData_authbusy;
  wire [1:0] DMINFORdData_authtype;
  wire [1:0] DMINFORdData_version;
  wire  HALTSUMRdData_serialfull;
  wire  HALTSUMRdData_serialvalid;
  wire [31:0] HALTSUMRdData_acks;
  wire  RAMWrData_interrupt;
  wire  RAMWrData_haltnot;
  wire [31:0] RAMWrData_data;
  wire  RAMRdData_interrupt;
  wire  RAMRdData_haltnot;
  wire [31:0] RAMRdData_data;
  wire  SETHALTNOTWrEn;
  wire [9:0] SETHALTNOTWrData;
  wire  CLEARDEBINTWrEn;
  wire [9:0] CLEARDEBINTWrData;
  wire  T_655_0;
  reg  interruptRegs_0;
  reg [31:0] GEN_111;
  wire  T_666_0;
  reg  haltnotRegs_0;
  reg [31:0] GEN_112;
  wire [31:0] haltnotStatus_0;
  wire [31:0] rdHaltnotStatus;
  wire [31:0] GEN_109;
  wire  haltnotSummary;
  reg [63:0] ramMem [0:7];
  reg [63:0] GEN_113;
  wire [63:0] ramMem_T_853_data;
  wire [2:0] ramMem_T_853_addr;
  wire  ramMem_T_853_en;
  wire [63:0] ramMem_T_854_data;
  wire [2:0] ramMem_T_854_addr;
  wire  ramMem_T_854_mask;
  wire  ramMem_T_854_en;
  wire [2:0] ramAddr;
  wire [63:0] ramRdData;
  wire [63:0] ramWrData;
  wire [63:0] ramWrMask;
  wire  ramWrEn;
  wire [3:0] dbRamAddr;
  wire [31:0] dbRamRdData;
  wire [31:0] dbRamWrData;
  wire  dbRamWrEn;
  wire  dbRamRdEn;
  wire [2:0] sbRamAddr;
  wire [63:0] sbRamRdData;
  wire [63:0] sbRamWrData;
  wire  sbRamWrEn;
  wire  sbRamRdEn;
  wire [63:0] sbRomRdData;
  wire  dbRdEn;
  wire  dbWrEn;
  wire [33:0] dbRdData;
  reg  dbStateReg;
  reg [31:0] GEN_122;
  wire [1:0] dbResult_resp;
  wire [33:0] dbResult_data;
  wire [4:0] dbReq_addr;
  wire [1:0] dbReq_op;
  wire [33:0] dbReq_data;
  reg [1:0] dbRespReg_resp;
  reg [31:0] GEN_123;
  reg [33:0] dbRespReg_data;
  reg [63:0] GEN_124;
  wire  rdCondWrFailure;
  wire  dbWrNeeded;
  wire [11:0] sbAddr;
  wire [63:0] sbRdData;
  wire [63:0] sbWrData;
  wire [63:0] sbWrMask;
  wire  sbWrEn;
  wire  sbRdEn;
  wire  stallFromDb;
  wire  stallFromSb;
  wire [9:0] GEN_110;
  wire  T_720;
  wire  T_721;
  wire  GEN_11;
  wire  GEN_12;
  wire  T_723;
  wire  T_724;
  wire  T_726;
  wire  T_727;
  wire  GEN_13;
  wire  GEN_14;
  wire  T_731;
  wire  T_732;
  wire  T_733;
  wire  T_735;
  wire  GEN_15;
  wire  GEN_16;
  wire  T_738;
  wire  GEN_17;
  wire  GEN_18;
  wire  T_741;
  wire  T_742;
  wire  T_745;
  wire  GEN_19;
  wire  GEN_20;
  wire  T_750;
  wire  T_751;
  wire  T_754;
  wire  GEN_21;
  wire  GEN_22;
  wire [3:0] T_782;
  wire [2:0] T_783;
  wire [31:0] T_801_0;
  wire [31:0] T_801_1;
  wire [31:0] dbRamWrMask_0;
  wire [31:0] dbRamWrMask_1;
  wire  T_806;
  wire [31:0] T_807;
  wire [31:0] T_808;
  wire [31:0] T_814_0;
  wire [31:0] T_814_1;
  wire [31:0] T_823_0;
  wire [31:0] T_823_1;
  wire [31:0] GEN_0;
  wire [31:0] GEN_23;
  wire [31:0] GEN_24;
  wire [31:0] GEN_1;
  wire [31:0] GEN_25;
  wire [63:0] T_831;
  wire [63:0] T_832;
  wire  T_833;
  wire  T_834;
  wire  T_835;
  wire  T_837;
  wire  T_838;
  wire  T_840;
  wire [63:0] dbRamWrDataVec;
  wire [63:0] T_841;
  wire [63:0] T_842;
  wire [63:0] T_843;
  wire [63:0] T_844;
  wire [63:0] T_845;
  wire [63:0] T_848;
  wire [63:0] T_849;
  wire  T_850;
  wire [2:0] T_851;
  wire [2:0] T_852;
  wire  T_855;
  wire  T_878_interrupt;
  wire  T_878_haltnot;
  wire [9:0] T_878_reserved0;
  wire [2:0] T_878_buserror;
  wire [2:0] T_878_serial;
  wire  T_878_autoincrement;
  wire [2:0] T_878_access;
  wire [9:0] T_878_hartid;
  wire  T_878_ndreset;
  wire  T_878_fullreset;
  wire  T_889;
  wire  T_890;
  wire [9:0] T_891;
  wire [2:0] T_892;
  wire  T_893;
  wire [2:0] T_894;
  wire [2:0] T_895;
  wire [9:0] T_896;
  wire  T_897;
  wire  T_898;
  wire  T_907_interrupt;
  wire  T_907_haltnot;
  wire [31:0] T_907_data;
  wire [31:0] T_911;
  wire  T_916;
  wire  T_918;
  wire  GEN_31;
  wire  T_920;
  wire  T_922;
  wire  T_923;
  wire  GEN_32;
  wire  T_927;
  wire  T_928;
  wire  GEN_33;
  wire  GEN_34;
  wire [9:0] GEN_35;
  wire [2:0] GEN_36;
  wire [2:0] GEN_37;
  wire  GEN_38;
  wire [2:0] GEN_39;
  wire [9:0] GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  T_931;
  wire  T_932;
  wire  T_933;
  wire  GEN_44;
  wire  T_936;
  wire  T_938;
  wire [1:0] T_941;
  wire  T_942;
  wire  T_943;
  wire  GEN_45;
  wire [9:0] GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  T_948;
  wire  GEN_49;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire [4:0] GEN_114;
  wire  T_961;
  wire [31:0] GEN_50;
  wire [1:0] T_966;
  wire [33:0] T_967;
  wire [33:0] GEN_51;
  wire [1:0] T_973;
  wire [3:0] T_974;
  wire [13:0] T_975;
  wire [15:0] T_976;
  wire [5:0] T_977;
  wire [1:0] T_978;
  wire [11:0] T_979;
  wire [17:0] T_980;
  wire [33:0] T_981;
  wire [33:0] GEN_53;
  wire  T_983;
  wire  T_989;
  wire [2:0] T_990;
  wire [4:0] T_991;
  wire [3:0] T_992;
  wire [6:0] T_993;
  wire [10:0] T_994;
  wire [15:0] T_995;
  wire [1:0] T_996;
  wire [1:0] T_997;
  wire [3:0] T_998;
  wire [4:0] T_999;
  wire [8:0] T_1000;
  wire [13:0] T_1001;
  wire [17:0] T_1002;
  wire [33:0] T_1003;
  wire [33:0] GEN_54;
  wire  T_1005;
  wire  T_1012;
  wire  T_1013;
  wire  T_1014;
  wire [33:0] GEN_55;
  wire [2:0] T_1016;
  wire  T_1018;
  wire  T_1028;
  wire  T_1029;
  wire  T_1030;
  wire [33:0] GEN_56;
  wire  T_1043;
  wire  T_1044;
  wire [33:0] GEN_57;
  wire  T_1046;
  wire  T_1048;
  wire  T_1049;
  wire  T_1051;
  wire  T_1054;
  wire  T_1055;
  wire  T_1056;
  wire [1:0] T_1059;
  wire  T_1061;
  wire  T_1062;
  wire  T_1064;
  wire  T_1065;
  wire  T_1066;
  wire  T_1067;
  wire  T_1069;
  wire  T_1071;
  wire  GEN_58;
  wire [1:0] GEN_59;
  wire [33:0] GEN_60;
  wire  GEN_61;
  wire [1:0] GEN_62;
  wire [33:0] GEN_63;
  wire  T_1076;
  wire  T_1077;
  wire  GEN_64;
  wire [1:0] GEN_65;
  wire [33:0] GEN_66;
  wire  T_1081;
  wire  T_1082;
  wire  GEN_67;
  wire  GEN_68;
  wire [1:0] GEN_69;
  wire [33:0] GEN_70;
  wire [63:0] T_1104_0;
  wire [63:0] T_1104_1;
  wire [63:0] T_1104_2;
  wire [63:0] T_1104_3;
  wire [63:0] T_1104_4;
  wire [63:0] T_1104_5;
  wire [63:0] T_1104_6;
  wire [63:0] T_1104_7;
  wire [63:0] T_1104_8;
  wire [63:0] T_1104_9;
  wire [63:0] T_1104_10;
  wire [63:0] T_1104_11;
  wire [63:0] T_1104_12;
  wire [63:0] T_1104_13;
  wire [63:0] T_1104_14;
  wire [3:0] T_1107;
  wire [3:0] T_1108;
  wire [63:0] GEN_6;
  wire [3:0] GEN_115;
  wire [63:0] GEN_71;
  wire [3:0] GEN_116;
  wire [63:0] GEN_72;
  wire [3:0] GEN_117;
  wire [63:0] GEN_73;
  wire [3:0] GEN_118;
  wire [63:0] GEN_74;
  wire [3:0] GEN_119;
  wire [63:0] GEN_75;
  wire [3:0] GEN_120;
  wire [63:0] GEN_76;
  wire [3:0] GEN_121;
  wire [63:0] GEN_77;
  wire [63:0] GEN_78;
  wire [63:0] GEN_79;
  wire [63:0] GEN_80;
  wire [63:0] GEN_81;
  wire [63:0] GEN_82;
  wire [63:0] GEN_83;
  wire [63:0] GEN_84;
  wire [31:0] T_1112;
  wire [31:0] T_1113;
  wire [31:0] T_1119_0;
  wire [31:0] T_1119_1;
  wire [31:0] T_1121;
  wire [31:0] T_1122;
  wire [31:0] T_1128_0;
  wire [31:0] T_1128_1;
  wire [31:0] GEN_7;
  wire [31:0] GEN_8;
  wire [3:0] T_1134;
  wire  T_1136;
  wire  GEN_87;
  wire [8:0] T_1137;
  wire  T_1140;
  wire [31:0] GEN_9;
  wire  T_1144;
  wire  T_1145;
  wire  T_1146;
  wire  T_1150;
  wire [31:0] GEN_10;
  wire  T_1154;
  wire  T_1155;
  wire  T_1156;
  wire [63:0] GEN_91;
  wire  GEN_92;
  wire  T_1165;
  wire  T_1168;
  wire  T_1169;
  wire  T_1171;
  wire  T_1172;
  wire [63:0] GEN_93;
  wire  T_1176;
  wire  T_1177;
  wire [63:0] GEN_94;
  reg [25:0] sbAcqReg_addr_block;
  reg [31:0] GEN_125;
  reg [1:0] sbAcqReg_client_xact_id;
  reg [31:0] GEN_136;
  reg [2:0] sbAcqReg_addr_beat;
  reg [31:0] GEN_137;
  reg  sbAcqReg_is_builtin_type;
  reg [31:0] GEN_138;
  reg [2:0] sbAcqReg_a_type;
  reg [31:0] GEN_139;
  reg [11:0] sbAcqReg_union;
  reg [31:0] GEN_140;
  reg [63:0] sbAcqReg_data;
  reg [63:0] GEN_141;
  reg  sbAcqValidReg;
  reg [31:0] GEN_142;
  wire  T_1206;
  wire  sbReg_get;
  wire  T_1207;
  wire  sbReg_getblk;
  wire  T_1208;
  wire  sbReg_put;
  wire  T_1209;
  wire  sbReg_putblk;
  wire  sbMultibeat;
  wire [2:0] GEN_126;
  wire [3:0] T_1211;
  wire [2:0] sbBeatInc1;
  wire  sbLast;
  wire [2:0] T_1213;
  wire [28:0] T_1214;
  wire [31:0] T_1215;
  wire  T_1216;
  wire  T_1217;
  wire  T_1218;
  wire  T_1219;
  wire  T_1221;
  wire  T_1222;
  wire [7:0] GEN_127;
  wire [8:0] T_1226;
  wire [7:0] T_1227;
  wire [7:0] T_1233_0;
  wire  T_1241;
  wire [7:0] T_1242;
  wire [7:0] T_1244;
  wire [7:0] T_1245;
  wire  T_1246;
  wire  T_1247;
  wire  T_1248;
  wire  T_1249;
  wire  T_1250;
  wire  T_1251;
  wire  T_1252;
  wire  T_1253;
  wire [7:0] GEN_128;
  wire [8:0] T_1255;
  wire [7:0] T_1256;
  wire [7:0] GEN_129;
  wire [8:0] T_1258;
  wire [7:0] T_1259;
  wire [7:0] GEN_130;
  wire [8:0] T_1261;
  wire [7:0] T_1262;
  wire [7:0] GEN_131;
  wire [8:0] T_1264;
  wire [7:0] T_1265;
  wire [7:0] GEN_132;
  wire [8:0] T_1267;
  wire [7:0] T_1268;
  wire [7:0] GEN_133;
  wire [8:0] T_1270;
  wire [7:0] T_1271;
  wire [7:0] GEN_134;
  wire [8:0] T_1273;
  wire [7:0] T_1274;
  wire [7:0] GEN_135;
  wire [8:0] T_1276;
  wire [7:0] T_1277;
  wire [7:0] T_1283_0;
  wire [7:0] T_1283_1;
  wire [7:0] T_1283_2;
  wire [7:0] T_1283_3;
  wire [7:0] T_1283_4;
  wire [7:0] T_1283_5;
  wire [7:0] T_1283_6;
  wire [7:0] T_1283_7;
  wire [15:0] T_1285;
  wire [15:0] T_1286;
  wire [31:0] T_1287;
  wire [15:0] T_1288;
  wire [15:0] T_1289;
  wire [31:0] T_1290;
  wire [63:0] T_1291;
  wire  T_1292;
  wire [25:0] GEN_95;
  wire [1:0] GEN_96;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire [2:0] GEN_99;
  wire [11:0] GEN_100;
  wire [63:0] GEN_101;
  wire  GEN_102;
  wire  T_1294;
  wire  T_1296;
  wire  T_1297;
  wire  GEN_103;
  wire [2:0] GEN_104;
  wire  GEN_105;
  wire  T_1300;
  wire  GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire  T_1318;
  wire [2:0] T_1319;
  wire  T_1320;
  wire [2:0] T_1321;
  wire  T_1322;
  wire [2:0] T_1323;
  wire  T_1324;
  wire [2:0] T_1325;
  wire  T_1326;
  wire [2:0] T_1327;
  wire  T_1328;
  wire [2:0] T_1329;
  wire  T_1330;
  wire [2:0] T_1331;
  wire [2:0] T_1355_addr_beat;
  wire [1:0] T_1355_client_xact_id;
  wire  T_1355_manager_xact_id;
  wire  T_1355_is_builtin_type;
  wire [3:0] T_1355_g_type;
  wire [63:0] T_1355_data;
  wire  T_1380;
  wire  T_1381;
  wire  T_1383;
  wire  T_1384;
  wire  T_1385;
  wire  sbStall;
  wire  T_1387;
  assign io_db_req_ready = T_1067;
  assign io_db_resp_valid = dbStateReg;
  assign io_db_resp_bits_resp = dbRespReg_resp;
  assign io_db_resp_bits_data = dbRespReg_data;
  assign io_debugInterrupts_0 = interruptRegs_0;
  assign io_tl_acquire_ready = T_1387;
  assign io_tl_grant_valid = sbAcqValidReg;
  assign io_tl_grant_bits_addr_beat = T_1355_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_1355_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_1355_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_1355_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_1355_g_type;
  assign io_tl_grant_bits_data = T_1355_data;
  assign io_ndreset = ndresetCtrReg;
  assign io_fullreset = CONTROLReg_fullreset;
  assign CONTROLReset_interrupt = 1'h0;
  assign CONTROLReset_haltnot = 1'h0;
  assign CONTROLReset_reserved0 = {{9'd0}, 1'h0};
  assign CONTROLReset_buserror = {{2'd0}, 1'h0};
  assign CONTROLReset_serial = {{2'd0}, 1'h0};
  assign CONTROLReset_autoincrement = 1'h0;
  assign CONTROLReset_access = {{1'd0}, 2'h2};
  assign CONTROLReset_hartid = {{9'd0}, 1'h0};
  assign CONTROLReset_ndreset = 1'h0;
  assign CONTROLReset_fullreset = 1'h0;
  assign CONTROLWrEn = GEN_32;
  assign CONTROLWrData_interrupt = T_878_interrupt;
  assign CONTROLWrData_haltnot = T_878_haltnot;
  assign CONTROLWrData_reserved0 = T_878_reserved0;
  assign CONTROLWrData_buserror = T_878_buserror;
  assign CONTROLWrData_serial = T_878_serial;
  assign CONTROLWrData_autoincrement = T_878_autoincrement;
  assign CONTROLWrData_access = T_878_access;
  assign CONTROLWrData_hartid = T_878_hartid;
  assign CONTROLWrData_ndreset = T_878_ndreset;
  assign CONTROLWrData_fullreset = T_878_fullreset;
  assign CONTROLRdData_interrupt = GEN_2;
  assign CONTROLRdData_haltnot = GEN_3;
  assign CONTROLRdData_reserved0 = CONTROLReg_reserved0;
  assign CONTROLRdData_buserror = CONTROLReg_buserror;
  assign CONTROLRdData_serial = CONTROLReg_serial;
  assign CONTROLRdData_autoincrement = CONTROLReg_autoincrement;
  assign CONTROLRdData_access = CONTROLReg_access;
  assign CONTROLRdData_hartid = CONTROLReg_hartid;
  assign CONTROLRdData_ndreset = ndresetCtrReg;
  assign CONTROLRdData_fullreset = CONTROLReg_fullreset;
  assign DMINFORdData_reserved0 = {{1'd0}, 1'h0};
  assign DMINFORdData_abussize = {{6'd0}, 1'h0};
  assign DMINFORdData_serialcount = {{3'd0}, 1'h0};
  assign DMINFORdData_access128 = 1'h0;
  assign DMINFORdData_access64 = 1'h0;
  assign DMINFORdData_access32 = 1'h0;
  assign DMINFORdData_access16 = 1'h0;
  assign DMINFORdData_accesss8 = 1'h0;
  assign DMINFORdData_dramsize = {{2'd0}, 4'hf};
  assign DMINFORdData_haltsum = 1'h0;
  assign DMINFORdData_reserved1 = {{2'd0}, 1'h0};
  assign DMINFORdData_authenticated = 1'h1;
  assign DMINFORdData_authbusy = 1'h0;
  assign DMINFORdData_authtype = {{1'd0}, 1'h0};
  assign DMINFORdData_version = {{1'd0}, 1'h1};
  assign HALTSUMRdData_serialfull = 1'h0;
  assign HALTSUMRdData_serialvalid = 1'h0;
  assign HALTSUMRdData_acks = {{31'd0}, haltnotSummary};
  assign RAMWrData_interrupt = T_907_interrupt;
  assign RAMWrData_haltnot = T_907_haltnot;
  assign RAMWrData_data = T_907_data;
  assign RAMRdData_interrupt = GEN_4;
  assign RAMRdData_haltnot = GEN_5;
  assign RAMRdData_data = dbRamRdData;
  assign SETHALTNOTWrEn = T_1146;
  assign SETHALTNOTWrData = GEN_7[9:0];
  assign CLEARDEBINTWrEn = T_1156;
  assign CLEARDEBINTWrData = GEN_8[9:0];
  assign T_655_0 = 1'h0;
  assign T_666_0 = 1'h0;
  assign haltnotStatus_0 = {{31'd0}, haltnotRegs_0};
  assign rdHaltnotStatus = GEN_50;
  assign GEN_109 = {{31'd0}, 1'h0};
  assign haltnotSummary = haltnotStatus_0 != GEN_109;
  assign ramMem_T_853_addr = ramAddr;
  assign ramMem_T_853_en = 1'h1;
  `ifdef SYNTHESIS
  assign ramMem_T_853_data = ramMem[ramMem_T_853_addr];
  `else
  assign ramMem_T_853_data = ramMem_T_853_addr >= 4'h8 ? $random : ramMem[ramMem_T_853_addr];
  `endif
  assign ramMem_T_854_data = ramWrData;
  assign ramMem_T_854_addr = ramAddr;
  assign ramMem_T_854_mask = ramWrEn;
  assign ramMem_T_854_en = ramWrEn;
  assign ramAddr = T_852;
  assign ramRdData = ramMem_T_853_data;
  assign ramWrData = T_849;
  assign ramWrMask = T_832;
  assign ramWrEn = T_855;
  assign dbRamAddr = T_782;
  assign dbRamRdData = GEN_1;
  assign dbRamWrData = dbReq_data[31:0];
  assign dbRamWrEn = GEN_31;
  assign dbRamRdEn = 1'h0;
  assign sbRamAddr = T_783;
  assign sbRamRdData = ramRdData;
  assign sbRamWrData = sbWrData;
  assign sbRamWrEn = GEN_87;
  assign sbRamRdEn = GEN_92;
  assign sbRomRdData = GEN_6;
  assign dbRdEn = T_1069;
  assign dbWrEn = T_1071;
  assign dbRdData = GEN_57;
  assign dbResult_resp = T_1059;
  assign dbResult_data = dbRdData;
  assign dbReq_addr = io_db_req_bits_addr;
  assign dbReq_op = io_db_req_bits_op;
  assign dbReq_data = io_db_req_bits_data;
  assign rdCondWrFailure = T_1049;
  assign dbWrNeeded = T_1056;
  assign sbAddr = T_1215[11:0];
  assign sbRdData = GEN_94;
  assign sbWrData = sbAcqReg_data;
  assign sbWrMask = T_1291;
  assign sbWrEn = T_1219;
  assign sbRdEn = T_1217;
  assign stallFromDb = 1'h0;
  assign stallFromSb = T_834;
  assign GEN_110 = {{9'd0}, 1'h0};
  assign T_720 = CONTROLWrData_hartid == GEN_110;
  assign T_721 = interruptRegs_0 | CONTROLWrData_interrupt;
  assign GEN_11 = T_720 ? T_721 : interruptRegs_0;
  assign GEN_12 = CONTROLWrEn ? GEN_11 : interruptRegs_0;
  assign T_723 = CONTROLWrEn == 1'h0;
  assign T_724 = T_723 & dbRamWrEn;
  assign T_726 = CONTROLReg_hartid == GEN_110;
  assign T_727 = interruptRegs_0 | RAMWrData_interrupt;
  assign GEN_13 = T_726 ? T_727 : GEN_12;
  assign GEN_14 = T_724 ? GEN_13 : GEN_12;
  assign T_731 = dbRamWrEn == 1'h0;
  assign T_732 = T_723 & T_731;
  assign T_733 = T_732 & CLEARDEBINTWrEn;
  assign T_735 = CLEARDEBINTWrData == 10'h0;
  assign GEN_15 = T_735 ? 1'h0 : GEN_14;
  assign GEN_16 = T_733 ? GEN_15 : GEN_14;
  assign T_738 = SETHALTNOTWrData == 10'h0;
  assign GEN_17 = T_738 ? 1'h1 : haltnotRegs_0;
  assign GEN_18 = SETHALTNOTWrEn ? GEN_17 : haltnotRegs_0;
  assign T_741 = SETHALTNOTWrEn == 1'h0;
  assign T_742 = T_741 & CONTROLWrEn;
  assign T_745 = haltnotRegs_0 & CONTROLWrData_haltnot;
  assign GEN_19 = T_720 ? T_745 : GEN_18;
  assign GEN_20 = T_742 ? GEN_19 : GEN_18;
  assign T_750 = T_741 & T_723;
  assign T_751 = T_750 & dbRamWrEn;
  assign T_754 = haltnotRegs_0 & RAMWrData_haltnot;
  assign GEN_21 = T_726 ? T_754 : GEN_20;
  assign GEN_22 = T_751 ? GEN_21 : GEN_20;
  assign T_782 = dbReq_addr[3:0];
  assign T_783 = sbAddr[5:3];
  assign T_801_0 = 32'hffffffff;
  assign T_801_1 = 32'hffffffff;
  assign dbRamWrMask_0 = GEN_23;
  assign dbRamWrMask_1 = GEN_24;
  assign T_806 = dbRamAddr[0];
  assign T_807 = ramRdData[31:0];
  assign T_808 = ramRdData[63:32];
  assign T_814_0 = T_807;
  assign T_814_1 = T_808;
  assign T_823_0 = 32'h0;
  assign T_823_1 = 32'h0;
  assign GEN_0 = 32'hffffffff;
  assign GEN_23 = 1'h0 == T_806 ? GEN_0 : T_823_0;
  assign GEN_24 = T_806 ? GEN_0 : T_823_1;
  assign GEN_1 = GEN_25;
  assign GEN_25 = T_806 ? T_814_1 : T_814_0;
  assign T_831 = {dbRamWrMask_1,dbRamWrMask_0};
  assign T_832 = sbRamWrEn ? sbWrMask : T_831;
  assign T_833 = dbRamWrEn | dbRamRdEn;
  assign T_834 = sbRamRdEn | sbRamWrEn;
  assign T_835 = T_833 & T_834;
  assign T_837 = T_835 == 1'h0;
  assign T_838 = T_837 | reset;
  assign T_840 = T_838 == 1'h0;
  assign dbRamWrDataVec = {dbRamWrData,dbRamWrData};
  assign T_841 = ramWrMask & sbRamWrData;
  assign T_842 = ~ ramWrMask;
  assign T_843 = T_842 & ramRdData;
  assign T_844 = T_841 | T_843;
  assign T_845 = ramWrMask & dbRamWrDataVec;
  assign T_848 = T_845 | T_843;
  assign T_849 = sbRamWrEn ? T_844 : T_848;
  assign T_850 = sbRamWrEn | sbRamRdEn;
  assign T_851 = dbRamAddr[3:1];
  assign T_852 = T_850 ? sbRamAddr : T_851;
  assign T_855 = sbRamWrEn | dbRamWrEn;
  assign T_878_interrupt = T_898;
  assign T_878_haltnot = T_897;
  assign T_878_reserved0 = T_896;
  assign T_878_buserror = T_895;
  assign T_878_serial = T_894;
  assign T_878_autoincrement = T_893;
  assign T_878_access = T_892;
  assign T_878_hartid = T_891;
  assign T_878_ndreset = T_890;
  assign T_878_fullreset = T_889;
  assign T_889 = dbReq_data[0];
  assign T_890 = dbReq_data[1];
  assign T_891 = dbReq_data[11:2];
  assign T_892 = dbReq_data[14:12];
  assign T_893 = dbReq_data[15];
  assign T_894 = dbReq_data[18:16];
  assign T_895 = dbReq_data[21:19];
  assign T_896 = dbReq_data[31:22];
  assign T_897 = dbReq_data[32];
  assign T_898 = dbReq_data[33];
  assign T_907_interrupt = T_898;
  assign T_907_haltnot = T_897;
  assign T_907_data = T_911;
  assign T_911 = dbReq_data[31:0];
  assign T_916 = dbReq_addr[4:4];
  assign T_918 = T_916 == 1'h0;
  assign GEN_31 = T_918 ? dbWrEn : 1'h0;
  assign T_920 = dbReq_addr == 5'h10;
  assign T_922 = T_918 == 1'h0;
  assign T_923 = T_922 & T_920;
  assign GEN_32 = T_923 ? dbWrEn : 1'h0;
  assign T_927 = T_920 == 1'h0;
  assign T_928 = T_922 & T_927;
  assign GEN_33 = reset ? CONTROLReset_interrupt : CONTROLReg_interrupt;
  assign GEN_34 = reset ? CONTROLReset_haltnot : CONTROLReg_haltnot;
  assign GEN_35 = reset ? CONTROLReset_reserved0 : CONTROLReg_reserved0;
  assign GEN_36 = reset ? CONTROLReset_buserror : CONTROLReg_buserror;
  assign GEN_37 = reset ? CONTROLReset_serial : CONTROLReg_serial;
  assign GEN_38 = reset ? CONTROLReset_autoincrement : CONTROLReg_autoincrement;
  assign GEN_39 = reset ? CONTROLReset_access : CONTROLReg_access;
  assign GEN_40 = reset ? CONTROLReset_hartid : CONTROLReg_hartid;
  assign GEN_41 = reset ? CONTROLReset_ndreset : CONTROLReg_ndreset;
  assign GEN_42 = reset ? CONTROLReset_fullreset : CONTROLReg_fullreset;
  assign GEN_43 = reset ? 1'h0 : ndresetCtrReg;
  assign T_931 = reset == 1'h0;
  assign T_932 = T_931 & CONTROLWrEn;
  assign T_933 = CONTROLReg_fullreset | CONTROLWrData_fullreset;
  assign GEN_44 = CONTROLWrData_ndreset ? 1'h1 : GEN_43;
  assign T_936 = CONTROLWrData_ndreset == 1'h0;
  assign T_938 = ndresetCtrReg == 1'h0;
  assign T_941 = ndresetCtrReg - 1'h1;
  assign T_942 = T_941[0:0];
  assign T_943 = T_938 ? 1'h0 : T_942;
  assign GEN_45 = T_936 ? T_943 : GEN_44;
  assign GEN_46 = T_932 ? CONTROLWrData_hartid : GEN_40;
  assign GEN_47 = T_932 ? T_933 : GEN_42;
  assign GEN_48 = T_932 ? GEN_45 : GEN_43;
  assign T_948 = T_931 & T_723;
  assign GEN_49 = T_948 ? T_943 : GEN_48;
  assign GEN_2 = interruptRegs_0;
  assign GEN_3 = haltnotRegs_0;
  assign GEN_4 = interruptRegs_0;
  assign GEN_5 = haltnotRegs_0;
  assign GEN_114 = {{4'd0}, 1'h0};
  assign T_961 = dbReq_addr == GEN_114;
  assign GEN_50 = T_961 ? haltnotStatus_0 : {{31'd0}, 1'h0};
  assign T_966 = {RAMRdData_interrupt,RAMRdData_haltnot};
  assign T_967 = {T_966,RAMRdData_data};
  assign GEN_51 = T_918 ? T_967 : {{33'd0}, 1'h0};
  assign T_973 = {CONTROLRdData_ndreset,CONTROLRdData_fullreset};
  assign T_974 = {CONTROLRdData_autoincrement,CONTROLRdData_access};
  assign T_975 = {T_974,CONTROLRdData_hartid};
  assign T_976 = {T_975,T_973};
  assign T_977 = {CONTROLRdData_buserror,CONTROLRdData_serial};
  assign T_978 = {CONTROLRdData_interrupt,CONTROLRdData_haltnot};
  assign T_979 = {T_978,CONTROLRdData_reserved0};
  assign T_980 = {T_979,T_977};
  assign T_981 = {T_980,T_976};
  assign GEN_53 = T_923 ? T_981 : GEN_51;
  assign T_983 = dbReq_addr == 5'h11;
  assign T_989 = T_928 & T_983;
  assign T_990 = {DMINFORdData_authbusy,DMINFORdData_authtype};
  assign T_991 = {T_990,DMINFORdData_version};
  assign T_992 = {DMINFORdData_reserved1,DMINFORdData_authenticated};
  assign T_993 = {DMINFORdData_dramsize,DMINFORdData_haltsum};
  assign T_994 = {T_993,T_992};
  assign T_995 = {T_994,T_991};
  assign T_996 = {DMINFORdData_access16,DMINFORdData_accesss8};
  assign T_997 = {DMINFORdData_access64,DMINFORdData_access32};
  assign T_998 = {T_997,T_996};
  assign T_999 = {DMINFORdData_serialcount,DMINFORdData_access128};
  assign T_1000 = {DMINFORdData_reserved0,DMINFORdData_abussize};
  assign T_1001 = {T_1000,T_999};
  assign T_1002 = {T_1001,T_998};
  assign T_1003 = {T_1002,T_995};
  assign GEN_54 = T_989 ? T_1003 : GEN_53;
  assign T_1005 = dbReq_addr == 5'h1b;
  assign T_1012 = T_983 == 1'h0;
  assign T_1013 = T_928 & T_1012;
  assign T_1014 = T_1013 & T_1005;
  assign GEN_55 = T_1014 ? {{33'd0}, 1'h0} : GEN_54;
  assign T_1016 = dbReq_addr[4:2];
  assign T_1018 = T_1016 == 3'h7;
  assign T_1028 = T_1005 == 1'h0;
  assign T_1029 = T_1013 & T_1028;
  assign T_1030 = T_1029 & T_1018;
  assign GEN_56 = T_1030 ? {{2'd0}, rdHaltnotStatus} : GEN_55;
  assign T_1043 = T_1018 == 1'h0;
  assign T_1044 = T_1029 & T_1043;
  assign GEN_57 = T_1044 ? {{33'd0}, 1'h0} : GEN_56;
  assign T_1046 = dbRdData[33];
  assign T_1048 = dbReq_op == 2'h3;
  assign T_1049 = T_1046 & T_1048;
  assign T_1051 = dbReq_op == 2'h2;
  assign T_1054 = ~ rdCondWrFailure;
  assign T_1055 = T_1048 & T_1054;
  assign T_1056 = T_1051 | T_1055;
  assign T_1059 = rdCondWrFailure ? 2'h1 : 2'h0;
  assign T_1061 = stallFromSb == 1'h0;
  assign T_1062 = dbStateReg == 1'h0;
  assign T_1064 = io_db_resp_ready & io_db_resp_valid;
  assign T_1065 = dbStateReg & T_1064;
  assign T_1066 = T_1062 | T_1065;
  assign T_1067 = T_1061 & T_1066;
  assign T_1069 = io_db_req_ready & io_db_req_valid;
  assign T_1071 = dbWrNeeded & T_1069;
  assign GEN_58 = T_1069 ? 1'h1 : dbStateReg;
  assign GEN_59 = T_1069 ? dbResult_resp : dbRespReg_resp;
  assign GEN_60 = T_1069 ? dbResult_data : dbRespReg_data;
  assign GEN_61 = T_1062 ? GEN_58 : dbStateReg;
  assign GEN_62 = T_1062 ? GEN_59 : dbRespReg_resp;
  assign GEN_63 = T_1062 ? GEN_60 : dbRespReg_data;
  assign T_1076 = T_1062 == 1'h0;
  assign T_1077 = T_1076 & dbStateReg;
  assign GEN_64 = T_1069 ? 1'h1 : GEN_61;
  assign GEN_65 = T_1069 ? dbResult_resp : GEN_62;
  assign GEN_66 = T_1069 ? dbResult_data : GEN_63;
  assign T_1081 = T_1069 == 1'h0;
  assign T_1082 = T_1081 & T_1064;
  assign GEN_67 = T_1082 ? 1'h0 : GEN_64;
  assign GEN_68 = T_1077 ? GEN_67 : GEN_61;
  assign GEN_69 = T_1077 ? GEN_65 : GEN_62;
  assign GEN_70 = T_1077 ? GEN_66 : GEN_63;
  assign T_1104_0 = 64'hc0006f03c0006f;
  assign T_1104_1 = 64'h80006ffff00413;
  assign T_1104_2 = 64'hff0000f00000413;
  assign T_1104_3 = 64'h42802e2343803483;
  assign T_1104_4 = 64'h10802023f1402473;
  assign T_1104_5 = 64'h8474137b002473;
  assign T_1104_6 = 64'h7b20247302041a63;
  assign T_1104_7 = 64'h7b2410737b200073;
  assign T_1104_8 = 64'h1c0474137b002473;
  assign T_1104_9 = 64'h41663f4040413;
  assign T_1104_10 = 64'h4000006742903c23;
  assign T_1104_11 = 64'h10802623f1402473;
  assign T_1104_12 = 64'h7b0024737b046073;
  assign T_1104_13 = 64'hfe040ce302047413;
  assign T_1104_14 = 64'hfe1ff06f;
  assign T_1107 = T_1108;
  assign T_1108 = sbAddr[6:3];
  assign GEN_6 = GEN_84;
  assign GEN_115 = {{3'd0}, 1'h1};
  assign GEN_71 = GEN_115 == T_1107 ? T_1104_1 : T_1104_0;
  assign GEN_116 = {{2'd0}, 2'h2};
  assign GEN_72 = GEN_116 == T_1107 ? T_1104_2 : GEN_71;
  assign GEN_117 = {{2'd0}, 2'h3};
  assign GEN_73 = GEN_117 == T_1107 ? T_1104_3 : GEN_72;
  assign GEN_118 = {{1'd0}, 3'h4};
  assign GEN_74 = GEN_118 == T_1107 ? T_1104_4 : GEN_73;
  assign GEN_119 = {{1'd0}, 3'h5};
  assign GEN_75 = GEN_119 == T_1107 ? T_1104_5 : GEN_74;
  assign GEN_120 = {{1'd0}, 3'h6};
  assign GEN_76 = GEN_120 == T_1107 ? T_1104_6 : GEN_75;
  assign GEN_121 = {{1'd0}, 3'h7};
  assign GEN_77 = GEN_121 == T_1107 ? T_1104_7 : GEN_76;
  assign GEN_78 = 4'h8 == T_1107 ? T_1104_8 : GEN_77;
  assign GEN_79 = 4'h9 == T_1107 ? T_1104_9 : GEN_78;
  assign GEN_80 = 4'ha == T_1107 ? T_1104_10 : GEN_79;
  assign GEN_81 = 4'hb == T_1107 ? T_1104_11 : GEN_80;
  assign GEN_82 = 4'hc == T_1107 ? T_1104_12 : GEN_81;
  assign GEN_83 = 4'hd == T_1107 ? T_1104_13 : GEN_82;
  assign GEN_84 = 4'he == T_1107 ? T_1104_14 : GEN_83;
  assign T_1112 = sbWrData[31:0];
  assign T_1113 = sbWrData[63:32];
  assign T_1119_0 = T_1112;
  assign T_1119_1 = T_1113;
  assign T_1121 = sbWrMask[31:0];
  assign T_1122 = sbWrMask[63:32];
  assign T_1128_0 = T_1121;
  assign T_1128_1 = T_1122;
  assign GEN_7 = T_1119_1;
  assign GEN_8 = T_1119_0;
  assign T_1134 = sbAddr[11:8];
  assign T_1136 = T_1134 == GEN_118;
  assign GEN_87 = T_1136 ? sbWrEn : 1'h0;
  assign T_1137 = sbAddr[11:3];
  assign T_1140 = T_1137 == 9'h21;
  assign GEN_9 = T_1128_1;
  assign T_1144 = GEN_9 != GEN_109;
  assign T_1145 = T_1140 & T_1144;
  assign T_1146 = T_1145 & sbWrEn;
  assign T_1150 = T_1137 == 9'h20;
  assign GEN_10 = T_1128_0;
  assign T_1154 = GEN_10 != GEN_109;
  assign T_1155 = T_1150 & T_1154;
  assign T_1156 = T_1155 & sbWrEn;
  assign GEN_91 = T_1136 ? sbRamRdData : {{63'd0}, 1'h0};
  assign GEN_92 = T_1136 ? sbRdEn : 1'h0;
  assign T_1165 = T_1134 == 4'h8;
  assign T_1168 = T_1134 == 4'h9;
  assign T_1169 = T_1165 | T_1168;
  assign T_1171 = T_1136 == 1'h0;
  assign T_1172 = T_1171 & T_1169;
  assign GEN_93 = T_1172 ? sbRomRdData : GEN_91;
  assign T_1176 = T_1169 == 1'h0;
  assign T_1177 = T_1171 & T_1176;
  assign GEN_94 = T_1177 ? {{63'd0}, 1'h0} : GEN_93;
  assign T_1206 = sbAcqReg_a_type == 3'h0;
  assign sbReg_get = sbAcqReg_is_builtin_type & T_1206;
  assign T_1207 = sbAcqReg_a_type == 3'h1;
  assign sbReg_getblk = sbAcqReg_is_builtin_type & T_1207;
  assign T_1208 = sbAcqReg_a_type == 3'h2;
  assign sbReg_put = sbAcqReg_is_builtin_type & T_1208;
  assign T_1209 = sbAcqReg_a_type == 3'h3;
  assign sbReg_putblk = sbAcqReg_is_builtin_type & T_1209;
  assign sbMultibeat = sbReg_getblk & sbAcqValidReg;
  assign GEN_126 = {{2'd0}, 1'h1};
  assign T_1211 = sbAcqReg_addr_beat + GEN_126;
  assign sbBeatInc1 = T_1211[2:0];
  assign sbLast = sbAcqReg_addr_beat == 3'h7;
  assign T_1213 = sbAcqReg_union[11:9];
  assign T_1214 = {sbAcqReg_addr_block,sbAcqReg_addr_beat};
  assign T_1215 = {T_1214,T_1213};
  assign T_1216 = sbReg_get | sbReg_getblk;
  assign T_1217 = sbAcqValidReg & T_1216;
  assign T_1218 = sbReg_put | sbReg_putblk;
  assign T_1219 = sbAcqValidReg & T_1218;
  assign T_1221 = sbAcqReg_a_type == 3'h4;
  assign T_1222 = sbAcqReg_is_builtin_type & T_1221;
  assign GEN_127 = {{7'd0}, 1'h1};
  assign T_1226 = 8'h0 - GEN_127;
  assign T_1227 = T_1226[7:0];
  assign T_1233_0 = T_1227;
  assign T_1241 = sbReg_putblk | sbReg_put;
  assign T_1242 = sbAcqReg_union[8:1];
  assign T_1244 = T_1241 ? T_1242 : {{7'd0}, 1'h0};
  assign T_1245 = T_1222 ? T_1233_0 : T_1244;
  assign T_1246 = T_1245[0];
  assign T_1247 = T_1245[1];
  assign T_1248 = T_1245[2];
  assign T_1249 = T_1245[3];
  assign T_1250 = T_1245[4];
  assign T_1251 = T_1245[5];
  assign T_1252 = T_1245[6];
  assign T_1253 = T_1245[7];
  assign GEN_128 = {{7'd0}, T_1246};
  assign T_1255 = 8'h0 - GEN_128;
  assign T_1256 = T_1255[7:0];
  assign GEN_129 = {{7'd0}, T_1247};
  assign T_1258 = 8'h0 - GEN_129;
  assign T_1259 = T_1258[7:0];
  assign GEN_130 = {{7'd0}, T_1248};
  assign T_1261 = 8'h0 - GEN_130;
  assign T_1262 = T_1261[7:0];
  assign GEN_131 = {{7'd0}, T_1249};
  assign T_1264 = 8'h0 - GEN_131;
  assign T_1265 = T_1264[7:0];
  assign GEN_132 = {{7'd0}, T_1250};
  assign T_1267 = 8'h0 - GEN_132;
  assign T_1268 = T_1267[7:0];
  assign GEN_133 = {{7'd0}, T_1251};
  assign T_1270 = 8'h0 - GEN_133;
  assign T_1271 = T_1270[7:0];
  assign GEN_134 = {{7'd0}, T_1252};
  assign T_1273 = 8'h0 - GEN_134;
  assign T_1274 = T_1273[7:0];
  assign GEN_135 = {{7'd0}, T_1253};
  assign T_1276 = 8'h0 - GEN_135;
  assign T_1277 = T_1276[7:0];
  assign T_1283_0 = T_1256;
  assign T_1283_1 = T_1259;
  assign T_1283_2 = T_1262;
  assign T_1283_3 = T_1265;
  assign T_1283_4 = T_1268;
  assign T_1283_5 = T_1271;
  assign T_1283_6 = T_1274;
  assign T_1283_7 = T_1277;
  assign T_1285 = {T_1283_1,T_1283_0};
  assign T_1286 = {T_1283_3,T_1283_2};
  assign T_1287 = {T_1286,T_1285};
  assign T_1288 = {T_1283_5,T_1283_4};
  assign T_1289 = {T_1283_7,T_1283_6};
  assign T_1290 = {T_1289,T_1288};
  assign T_1291 = {T_1290,T_1287};
  assign T_1292 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign GEN_95 = T_1292 ? io_tl_acquire_bits_addr_block : sbAcqReg_addr_block;
  assign GEN_96 = T_1292 ? io_tl_acquire_bits_client_xact_id : sbAcqReg_client_xact_id;
  assign GEN_97 = T_1292 ? io_tl_acquire_bits_addr_beat : sbAcqReg_addr_beat;
  assign GEN_98 = T_1292 ? io_tl_acquire_bits_is_builtin_type : sbAcqReg_is_builtin_type;
  assign GEN_99 = T_1292 ? io_tl_acquire_bits_a_type : sbAcqReg_a_type;
  assign GEN_100 = T_1292 ? io_tl_acquire_bits_union : sbAcqReg_union;
  assign GEN_101 = T_1292 ? io_tl_acquire_bits_data : sbAcqReg_data;
  assign GEN_102 = T_1292 ? 1'h1 : sbAcqValidReg;
  assign T_1294 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_1296 = T_1292 == 1'h0;
  assign T_1297 = T_1296 & T_1294;
  assign GEN_103 = sbLast ? 1'h0 : GEN_102;
  assign GEN_104 = sbMultibeat ? sbBeatInc1 : GEN_97;
  assign GEN_105 = sbMultibeat ? GEN_103 : GEN_102;
  assign T_1300 = sbMultibeat == 1'h0;
  assign GEN_106 = T_1300 ? 1'h0 : GEN_105;
  assign GEN_107 = T_1297 ? GEN_104 : GEN_97;
  assign GEN_108 = T_1297 ? GEN_106 : GEN_102;
  assign T_1318 = 3'h6 == sbAcqReg_a_type;
  assign T_1319 = T_1318 ? 3'h1 : 3'h3;
  assign T_1320 = 3'h5 == sbAcqReg_a_type;
  assign T_1321 = T_1320 ? 3'h1 : T_1319;
  assign T_1322 = 3'h4 == sbAcqReg_a_type;
  assign T_1323 = T_1322 ? 3'h4 : T_1321;
  assign T_1324 = 3'h3 == sbAcqReg_a_type;
  assign T_1325 = T_1324 ? 3'h3 : T_1323;
  assign T_1326 = 3'h2 == sbAcqReg_a_type;
  assign T_1327 = T_1326 ? 3'h3 : T_1325;
  assign T_1328 = 3'h1 == sbAcqReg_a_type;
  assign T_1329 = T_1328 ? 3'h5 : T_1327;
  assign T_1330 = 3'h0 == sbAcqReg_a_type;
  assign T_1331 = T_1330 ? 3'h4 : T_1329;
  assign T_1355_addr_beat = sbAcqReg_addr_beat;
  assign T_1355_client_xact_id = sbAcqReg_client_xact_id;
  assign T_1355_manager_xact_id = 1'h0;
  assign T_1355_is_builtin_type = 1'h1;
  assign T_1355_g_type = {{1'd0}, T_1331};
  assign T_1355_data = sbRdData;
  assign T_1380 = sbLast == 1'h0;
  assign T_1381 = sbMultibeat & T_1380;
  assign T_1383 = io_tl_grant_ready == 1'h0;
  assign T_1384 = io_tl_grant_valid & T_1383;
  assign T_1385 = T_1381 | T_1384;
  assign sbStall = T_1385 | stallFromDb;
  assign T_1387 = sbStall == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_26 = {1{$random}};
  CONTROLReg_interrupt = GEN_26[0:0];
  GEN_27 = {1{$random}};
  CONTROLReg_haltnot = GEN_27[0:0];
  GEN_28 = {1{$random}};
  CONTROLReg_reserved0 = GEN_28[9:0];
  GEN_29 = {1{$random}};
  CONTROLReg_buserror = GEN_29[2:0];
  GEN_30 = {1{$random}};
  CONTROLReg_serial = GEN_30[2:0];
  GEN_52 = {1{$random}};
  CONTROLReg_autoincrement = GEN_52[0:0];
  GEN_85 = {1{$random}};
  CONTROLReg_access = GEN_85[2:0];
  GEN_86 = {1{$random}};
  CONTROLReg_hartid = GEN_86[9:0];
  GEN_88 = {1{$random}};
  CONTROLReg_ndreset = GEN_88[0:0];
  GEN_89 = {1{$random}};
  CONTROLReg_fullreset = GEN_89[0:0];
  GEN_90 = {1{$random}};
  ndresetCtrReg = GEN_90[0:0];
  GEN_111 = {1{$random}};
  interruptRegs_0 = GEN_111[0:0];
  GEN_112 = {1{$random}};
  haltnotRegs_0 = GEN_112[0:0];
  GEN_113 = {2{$random}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ramMem[initvar] = GEN_113[63:0];
  GEN_122 = {1{$random}};
  dbStateReg = GEN_122[0:0];
  GEN_123 = {1{$random}};
  dbRespReg_resp = GEN_123[1:0];
  GEN_124 = {2{$random}};
  dbRespReg_data = GEN_124[33:0];
  GEN_125 = {1{$random}};
  sbAcqReg_addr_block = GEN_125[25:0];
  GEN_136 = {1{$random}};
  sbAcqReg_client_xact_id = GEN_136[1:0];
  GEN_137 = {1{$random}};
  sbAcqReg_addr_beat = GEN_137[2:0];
  GEN_138 = {1{$random}};
  sbAcqReg_is_builtin_type = GEN_138[0:0];
  GEN_139 = {1{$random}};
  sbAcqReg_a_type = GEN_139[2:0];
  GEN_140 = {1{$random}};
  sbAcqReg_union = GEN_140[11:0];
  GEN_141 = {2{$random}};
  sbAcqReg_data = GEN_141[63:0];
  GEN_142 = {1{$random}};
  sbAcqValidReg = GEN_142[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_interrupt <= CONTROLReset_interrupt;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_haltnot <= CONTROLReset_haltnot;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_reserved0 <= CONTROLReset_reserved0;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_buserror <= CONTROLReset_buserror;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_serial <= CONTROLReset_serial;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_autoincrement <= CONTROLReset_autoincrement;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_access <= CONTROLReset_access;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_932) begin
        CONTROLReg_hartid <= CONTROLWrData_hartid;
      end else begin
        if(reset) begin
          CONTROLReg_hartid <= CONTROLReset_hartid;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_ndreset <= CONTROLReset_ndreset;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_932) begin
        CONTROLReg_fullreset <= T_933;
      end else begin
        if(reset) begin
          CONTROLReg_fullreset <= CONTROLReset_fullreset;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_948) begin
        if(T_938) begin
          ndresetCtrReg <= 1'h0;
        end else begin
          ndresetCtrReg <= T_942;
        end
      end else begin
        if(T_932) begin
          if(T_936) begin
            if(T_938) begin
              ndresetCtrReg <= 1'h0;
            end else begin
              ndresetCtrReg <= T_942;
            end
          end else begin
            if(CONTROLWrData_ndreset) begin
              ndresetCtrReg <= 1'h1;
            end else begin
              if(reset) begin
                ndresetCtrReg <= 1'h0;
              end
            end
          end
        end else begin
          if(reset) begin
            ndresetCtrReg <= 1'h0;
          end
        end
      end
    end
    if(reset) begin
      interruptRegs_0 <= T_655_0;
    end else begin
      if(T_733) begin
        if(T_735) begin
          interruptRegs_0 <= 1'h0;
        end else begin
          if(T_724) begin
            if(T_726) begin
              interruptRegs_0 <= T_727;
            end else begin
              if(CONTROLWrEn) begin
                if(T_720) begin
                  interruptRegs_0 <= T_721;
                end
              end
            end
          end else begin
            if(CONTROLWrEn) begin
              if(T_720) begin
                interruptRegs_0 <= T_721;
              end
            end
          end
        end
      end else begin
        if(T_724) begin
          if(T_726) begin
            interruptRegs_0 <= T_727;
          end else begin
            if(CONTROLWrEn) begin
              if(T_720) begin
                interruptRegs_0 <= T_721;
              end
            end
          end
        end else begin
          if(CONTROLWrEn) begin
            if(T_720) begin
              interruptRegs_0 <= T_721;
            end
          end
        end
      end
    end
    if(reset) begin
      haltnotRegs_0 <= T_666_0;
    end else begin
      if(T_751) begin
        if(T_726) begin
          haltnotRegs_0 <= T_754;
        end else begin
          if(T_742) begin
            if(T_720) begin
              haltnotRegs_0 <= T_745;
            end else begin
              if(SETHALTNOTWrEn) begin
                if(T_738) begin
                  haltnotRegs_0 <= 1'h1;
                end
              end
            end
          end else begin
            if(SETHALTNOTWrEn) begin
              if(T_738) begin
                haltnotRegs_0 <= 1'h1;
              end
            end
          end
        end
      end else begin
        if(T_742) begin
          if(T_720) begin
            haltnotRegs_0 <= T_745;
          end else begin
            if(SETHALTNOTWrEn) begin
              if(T_738) begin
                haltnotRegs_0 <= 1'h1;
              end
            end
          end
        end else begin
          if(SETHALTNOTWrEn) begin
            if(T_738) begin
              haltnotRegs_0 <= 1'h1;
            end
          end
        end
      end
    end
    if(ramMem_T_854_en & ramMem_T_854_mask) begin
      ramMem[ramMem_T_854_addr] <= ramMem_T_854_data;
    end
    if(reset) begin
      dbStateReg <= 1'h0;
    end else begin
      if(T_1077) begin
        if(T_1082) begin
          dbStateReg <= 1'h0;
        end else begin
          if(T_1069) begin
            dbStateReg <= 1'h1;
          end else begin
            if(T_1062) begin
              if(T_1069) begin
                dbStateReg <= 1'h1;
              end
            end
          end
        end
      end else begin
        if(T_1062) begin
          if(T_1069) begin
            dbStateReg <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1077) begin
        if(T_1069) begin
          dbRespReg_resp <= dbResult_resp;
        end else begin
          if(T_1062) begin
            if(T_1069) begin
              dbRespReg_resp <= dbResult_resp;
            end
          end
        end
      end else begin
        if(T_1062) begin
          if(T_1069) begin
            dbRespReg_resp <= dbResult_resp;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1077) begin
        if(T_1069) begin
          dbRespReg_data <= dbResult_data;
        end else begin
          if(T_1062) begin
            if(T_1069) begin
              dbRespReg_data <= dbResult_data;
            end
          end
        end
      end else begin
        if(T_1062) begin
          if(T_1069) begin
            dbRespReg_data <= dbResult_data;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1292) begin
        sbAcqReg_addr_block <= io_tl_acquire_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1292) begin
        sbAcqReg_client_xact_id <= io_tl_acquire_bits_client_xact_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1297) begin
        if(sbMultibeat) begin
          sbAcqReg_addr_beat <= sbBeatInc1;
        end else begin
          if(T_1292) begin
            sbAcqReg_addr_beat <= io_tl_acquire_bits_addr_beat;
          end
        end
      end else begin
        if(T_1292) begin
          sbAcqReg_addr_beat <= io_tl_acquire_bits_addr_beat;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1292) begin
        sbAcqReg_is_builtin_type <= io_tl_acquire_bits_is_builtin_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1292) begin
        sbAcqReg_a_type <= io_tl_acquire_bits_a_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1292) begin
        sbAcqReg_union <= io_tl_acquire_bits_union;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1292) begin
        sbAcqReg_data <= io_tl_acquire_bits_data;
      end
    end
    if(reset) begin
      sbAcqValidReg <= 1'h0;
    end else begin
      if(T_1297) begin
        if(T_1300) begin
          sbAcqValidReg <= 1'h0;
        end else begin
          if(sbMultibeat) begin
            if(sbLast) begin
              sbAcqValidReg <= 1'h0;
            end else begin
              if(T_1292) begin
                sbAcqValidReg <= 1'h1;
              end
            end
          end else begin
            if(T_1292) begin
              sbAcqValidReg <= 1'h1;
            end
          end
        end
      end else begin
        if(T_1292) begin
          sbAcqValidReg <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_840) begin
          $fwrite(32'h80000002,"Assertion failed: Stall logic should have prevented concurrent SB/DB RAM Access\n    at Debug.scala:652 assert (!((dbRamWrEn | dbRamRdEn) & (sbRamRdEn | sbRamWrEn)), \"Stall logic should have prevented concurrent SB/DB RAM Access\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_840) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_840) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module PRCI(
  input   clk,
  input   reset,
  input   io_interrupts_0_meip,
  input   io_interrupts_0_seip,
  input   io_interrupts_0_debug,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_tiles_0_reset,
  output  io_tiles_0_id,
  output  io_tiles_0_interrupts_meip,
  output  io_tiles_0_interrupts_seip,
  output  io_tiles_0_interrupts_debug,
  output  io_tiles_0_interrupts_mtip,
  output  io_tiles_0_interrupts_msip,
  input   io_rtcTick
);
  reg [63:0] timecmp_0;
  reg [63:0] GEN_4;
  reg [63:0] time$;
  reg [63:0] GEN_5;
  wire [63:0] GEN_45;
  wire [64:0] T_525;
  wire [63:0] T_526;
  wire [63:0] GEN_0;
  wire [31:0] T_533_0;
  reg [31:0] ipi_0;
  reg [31:0] GEN_6;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire [2:0] T_561;
  wire [28:0] T_562;
  wire [31:0] T_563;
  wire [15:0] addr;
  wire [63:0] rdata;
  wire  T_583;
  wire [2:0] T_584;
  wire  T_585;
  wire [2:0] T_586;
  wire  T_587;
  wire [2:0] T_588;
  wire  T_589;
  wire [2:0] T_590;
  wire  T_591;
  wire [2:0] T_592;
  wire  T_593;
  wire [2:0] T_594;
  wire  T_595;
  wire [2:0] T_596;
  wire [2:0] T_621_addr_beat;
  wire [1:0] T_621_client_xact_id;
  wire  T_621_manager_xact_id;
  wire  T_621_is_builtin_type;
  wire [3:0] T_621_g_type;
  wire [63:0] T_621_data;
  wire  T_643;
  wire [63:0] GEN_46;
  wire [64:0] T_645;
  wire [63:0] T_646;
  wire [63:0] T_652_0;
  wire [63:0] GEN_2;
  wire [15:0] GEN_47;
  wire  T_658;
  wire  T_660;
  wire  T_661;
  wire  T_669;
  wire  T_670;
  wire [7:0] GEN_48;
  wire [8:0] T_674;
  wire [7:0] T_675;
  wire [7:0] T_681_0;
  wire  T_684;
  wire  T_685;
  wire  T_687;
  wire  T_688;
  wire  T_689;
  wire [7:0] T_690;
  wire [7:0] T_692;
  wire [7:0] T_693;
  wire  T_694;
  wire  T_695;
  wire  T_696;
  wire  T_697;
  wire  T_698;
  wire  T_699;
  wire  T_700;
  wire  T_701;
  wire [7:0] GEN_49;
  wire [8:0] T_703;
  wire [7:0] T_704;
  wire [7:0] GEN_50;
  wire [8:0] T_706;
  wire [7:0] T_707;
  wire [7:0] GEN_51;
  wire [8:0] T_709;
  wire [7:0] T_710;
  wire [7:0] GEN_52;
  wire [8:0] T_712;
  wire [7:0] T_713;
  wire [7:0] GEN_53;
  wire [8:0] T_715;
  wire [7:0] T_716;
  wire [7:0] GEN_54;
  wire [8:0] T_718;
  wire [7:0] T_719;
  wire [7:0] GEN_55;
  wire [8:0] T_721;
  wire [7:0] T_722;
  wire [7:0] GEN_56;
  wire [8:0] T_724;
  wire [7:0] T_725;
  wire [7:0] T_731_0;
  wire [7:0] T_731_1;
  wire [7:0] T_731_2;
  wire [7:0] T_731_3;
  wire [7:0] T_731_4;
  wire [7:0] T_731_5;
  wire [7:0] T_731_6;
  wire [7:0] T_731_7;
  wire [15:0] T_733;
  wire [15:0] T_734;
  wire [31:0] T_735;
  wire [15:0] T_736;
  wire [15:0] T_737;
  wire [31:0] T_738;
  wire [63:0] T_739;
  wire [63:0] T_740;
  wire [7:0] T_754_0;
  wire [7:0] T_766;
  wire  T_767;
  wire  T_768;
  wire  T_769;
  wire  T_770;
  wire  T_771;
  wire  T_772;
  wire  T_773;
  wire  T_774;
  wire [7:0] GEN_58;
  wire [8:0] T_776;
  wire [7:0] T_777;
  wire [7:0] GEN_59;
  wire [8:0] T_779;
  wire [7:0] T_780;
  wire [7:0] GEN_60;
  wire [8:0] T_782;
  wire [7:0] T_783;
  wire [7:0] GEN_61;
  wire [8:0] T_785;
  wire [7:0] T_786;
  wire [7:0] GEN_62;
  wire [8:0] T_788;
  wire [7:0] T_789;
  wire [7:0] GEN_63;
  wire [8:0] T_791;
  wire [7:0] T_792;
  wire [7:0] GEN_64;
  wire [8:0] T_794;
  wire [7:0] T_795;
  wire [7:0] GEN_65;
  wire [8:0] T_797;
  wire [7:0] T_798;
  wire [7:0] T_804_0;
  wire [7:0] T_804_1;
  wire [7:0] T_804_2;
  wire [7:0] T_804_3;
  wire [7:0] T_804_4;
  wire [7:0] T_804_5;
  wire [7:0] T_804_6;
  wire [7:0] T_804_7;
  wire [15:0] T_806;
  wire [15:0] T_807;
  wire [31:0] T_808;
  wire [15:0] T_809;
  wire [15:0] T_810;
  wire [31:0] T_811;
  wire [63:0] T_812;
  wire [63:0] T_813;
  wire [63:0] T_814;
  wire [63:0] T_815;
  wire [63:0] GEN_3;
  wire [63:0] GEN_22;
  wire [63:0] GEN_23;
  wire  T_827;
  wire  T_828;
  wire [7:0] T_848_0;
  wire [7:0] T_860;
  wire  T_861;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire  T_865;
  wire  T_866;
  wire  T_867;
  wire  T_868;
  wire [7:0] GEN_67;
  wire [8:0] T_870;
  wire [7:0] T_871;
  wire [7:0] GEN_68;
  wire [8:0] T_873;
  wire [7:0] T_874;
  wire [7:0] GEN_69;
  wire [8:0] T_876;
  wire [7:0] T_877;
  wire [7:0] GEN_70;
  wire [8:0] T_879;
  wire [7:0] T_880;
  wire [7:0] GEN_71;
  wire [8:0] T_882;
  wire [7:0] T_883;
  wire [7:0] GEN_72;
  wire [8:0] T_885;
  wire [7:0] T_886;
  wire [7:0] GEN_73;
  wire [8:0] T_888;
  wire [7:0] T_889;
  wire [7:0] GEN_74;
  wire [8:0] T_891;
  wire [7:0] T_892;
  wire [7:0] T_898_0;
  wire [7:0] T_898_1;
  wire [7:0] T_898_2;
  wire [7:0] T_898_3;
  wire [7:0] T_898_4;
  wire [7:0] T_898_5;
  wire [7:0] T_898_6;
  wire [7:0] T_898_7;
  wire [15:0] T_900;
  wire [15:0] T_901;
  wire [31:0] T_902;
  wire [15:0] T_903;
  wire [15:0] T_904;
  wire [31:0] T_905;
  wire [63:0] T_906;
  wire [63:0] T_907;
  wire [7:0] T_921_0;
  wire [7:0] T_933;
  wire  T_934;
  wire  T_935;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire  T_940;
  wire  T_941;
  wire [7:0] GEN_76;
  wire [8:0] T_943;
  wire [7:0] T_944;
  wire [7:0] GEN_77;
  wire [8:0] T_946;
  wire [7:0] T_947;
  wire [7:0] GEN_78;
  wire [8:0] T_949;
  wire [7:0] T_950;
  wire [7:0] GEN_79;
  wire [8:0] T_952;
  wire [7:0] T_953;
  wire [7:0] GEN_80;
  wire [8:0] T_955;
  wire [7:0] T_956;
  wire [7:0] GEN_81;
  wire [8:0] T_958;
  wire [7:0] T_959;
  wire [7:0] GEN_82;
  wire [8:0] T_961;
  wire [7:0] T_962;
  wire [7:0] GEN_83;
  wire [8:0] T_964;
  wire [7:0] T_965;
  wire [7:0] T_971_0;
  wire [7:0] T_971_1;
  wire [7:0] T_971_2;
  wire [7:0] T_971_3;
  wire [7:0] T_971_4;
  wire [7:0] T_971_5;
  wire [7:0] T_971_6;
  wire [7:0] T_971_7;
  wire [15:0] T_973;
  wire [15:0] T_974;
  wire [31:0] T_975;
  wire [15:0] T_976;
  wire [15:0] T_977;
  wire [31:0] T_978;
  wire [63:0] T_979;
  wire [63:0] T_980;
  wire [63:0] GEN_84;
  wire [63:0] T_981;
  wire [63:0] T_982;
  wire [63:0] GEN_24;
  wire [63:0] T_993;
  wire [63:0] GEN_43;
  wire [63:0] GEN_44;
  wire  T_994;
  wire  T_995;
  reg  GEN_1;
  reg [31:0] GEN_7;
  Queue_20 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_621_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_621_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_621_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_621_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_621_g_type;
  assign io_tl_grant_bits_data = T_621_data;
  assign io_tiles_0_reset = GEN_1;
  assign io_tiles_0_id = 1'h0;
  assign io_tiles_0_interrupts_meip = io_interrupts_0_meip;
  assign io_tiles_0_interrupts_seip = io_interrupts_0_seip;
  assign io_tiles_0_interrupts_debug = io_interrupts_0_debug;
  assign io_tiles_0_interrupts_mtip = T_995;
  assign io_tiles_0_interrupts_msip = T_994;
  assign GEN_45 = {{63'd0}, 1'h1};
  assign T_525 = time$ + GEN_45;
  assign T_526 = T_525[63:0];
  assign GEN_0 = io_rtcTick ? T_526 : time$;
  assign T_533_0 = 32'h0;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_561 = acq_io_deq_bits_union[11:9];
  assign T_562 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_563 = {T_562,T_561};
  assign addr = T_563[15:0];
  assign rdata = GEN_44;
  assign T_583 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_584 = T_583 ? 3'h1 : 3'h3;
  assign T_585 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_586 = T_585 ? 3'h1 : T_584;
  assign T_587 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_588 = T_587 ? 3'h4 : T_586;
  assign T_589 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_590 = T_589 ? 3'h3 : T_588;
  assign T_591 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_592 = T_591 ? 3'h3 : T_590;
  assign T_593 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_594 = T_593 ? 3'h5 : T_592;
  assign T_595 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_596 = T_595 ? 3'h4 : T_594;
  assign T_621_addr_beat = {{2'd0}, 1'h0};
  assign T_621_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_621_manager_xact_id = 1'h0;
  assign T_621_is_builtin_type = 1'h1;
  assign T_621_g_type = {{1'd0}, T_596};
  assign T_621_data = rdata;
  assign T_643 = addr[15];
  assign GEN_46 = {{63'd0}, 1'h0};
  assign T_645 = time$ + GEN_46;
  assign T_646 = T_645[63:0];
  assign T_652_0 = T_646;
  assign GEN_2 = T_643 ? T_652_0 : {{63'd0}, 1'h0};
  assign GEN_47 = {{1'd0}, 15'h4000};
  assign T_658 = addr >= GEN_47;
  assign T_660 = T_643 == 1'h0;
  assign T_661 = T_660 & T_658;
  assign T_669 = acq_io_deq_bits_a_type == 3'h4;
  assign T_670 = acq_io_deq_bits_is_builtin_type & T_669;
  assign GEN_48 = {{7'd0}, 1'h1};
  assign T_674 = 8'h0 - GEN_48;
  assign T_675 = T_674[7:0];
  assign T_681_0 = T_675;
  assign T_684 = acq_io_deq_bits_a_type == 3'h3;
  assign T_685 = acq_io_deq_bits_is_builtin_type & T_684;
  assign T_687 = acq_io_deq_bits_a_type == 3'h2;
  assign T_688 = acq_io_deq_bits_is_builtin_type & T_687;
  assign T_689 = T_685 | T_688;
  assign T_690 = acq_io_deq_bits_union[8:1];
  assign T_692 = T_689 ? T_690 : {{7'd0}, 1'h0};
  assign T_693 = T_670 ? T_681_0 : T_692;
  assign T_694 = T_693[0];
  assign T_695 = T_693[1];
  assign T_696 = T_693[2];
  assign T_697 = T_693[3];
  assign T_698 = T_693[4];
  assign T_699 = T_693[5];
  assign T_700 = T_693[6];
  assign T_701 = T_693[7];
  assign GEN_49 = {{7'd0}, T_694};
  assign T_703 = 8'h0 - GEN_49;
  assign T_704 = T_703[7:0];
  assign GEN_50 = {{7'd0}, T_695};
  assign T_706 = 8'h0 - GEN_50;
  assign T_707 = T_706[7:0];
  assign GEN_51 = {{7'd0}, T_696};
  assign T_709 = 8'h0 - GEN_51;
  assign T_710 = T_709[7:0];
  assign GEN_52 = {{7'd0}, T_697};
  assign T_712 = 8'h0 - GEN_52;
  assign T_713 = T_712[7:0];
  assign GEN_53 = {{7'd0}, T_698};
  assign T_715 = 8'h0 - GEN_53;
  assign T_716 = T_715[7:0];
  assign GEN_54 = {{7'd0}, T_699};
  assign T_718 = 8'h0 - GEN_54;
  assign T_719 = T_718[7:0];
  assign GEN_55 = {{7'd0}, T_700};
  assign T_721 = 8'h0 - GEN_55;
  assign T_722 = T_721[7:0];
  assign GEN_56 = {{7'd0}, T_701};
  assign T_724 = 8'h0 - GEN_56;
  assign T_725 = T_724[7:0];
  assign T_731_0 = T_704;
  assign T_731_1 = T_707;
  assign T_731_2 = T_710;
  assign T_731_3 = T_713;
  assign T_731_4 = T_716;
  assign T_731_5 = T_719;
  assign T_731_6 = T_722;
  assign T_731_7 = T_725;
  assign T_733 = {T_731_1,T_731_0};
  assign T_734 = {T_731_3,T_731_2};
  assign T_735 = {T_734,T_733};
  assign T_736 = {T_731_5,T_731_4};
  assign T_737 = {T_731_7,T_731_6};
  assign T_738 = {T_737,T_736};
  assign T_739 = {T_738,T_735};
  assign T_740 = acq_io_deq_bits_data & T_739;
  assign T_754_0 = T_675;
  assign T_766 = T_670 ? T_754_0 : T_692;
  assign T_767 = T_766[0];
  assign T_768 = T_766[1];
  assign T_769 = T_766[2];
  assign T_770 = T_766[3];
  assign T_771 = T_766[4];
  assign T_772 = T_766[5];
  assign T_773 = T_766[6];
  assign T_774 = T_766[7];
  assign GEN_58 = {{7'd0}, T_767};
  assign T_776 = 8'h0 - GEN_58;
  assign T_777 = T_776[7:0];
  assign GEN_59 = {{7'd0}, T_768};
  assign T_779 = 8'h0 - GEN_59;
  assign T_780 = T_779[7:0];
  assign GEN_60 = {{7'd0}, T_769};
  assign T_782 = 8'h0 - GEN_60;
  assign T_783 = T_782[7:0];
  assign GEN_61 = {{7'd0}, T_770};
  assign T_785 = 8'h0 - GEN_61;
  assign T_786 = T_785[7:0];
  assign GEN_62 = {{7'd0}, T_771};
  assign T_788 = 8'h0 - GEN_62;
  assign T_789 = T_788[7:0];
  assign GEN_63 = {{7'd0}, T_772};
  assign T_791 = 8'h0 - GEN_63;
  assign T_792 = T_791[7:0];
  assign GEN_64 = {{7'd0}, T_773};
  assign T_794 = 8'h0 - GEN_64;
  assign T_795 = T_794[7:0];
  assign GEN_65 = {{7'd0}, T_774};
  assign T_797 = 8'h0 - GEN_65;
  assign T_798 = T_797[7:0];
  assign T_804_0 = T_777;
  assign T_804_1 = T_780;
  assign T_804_2 = T_783;
  assign T_804_3 = T_786;
  assign T_804_4 = T_789;
  assign T_804_5 = T_792;
  assign T_804_6 = T_795;
  assign T_804_7 = T_798;
  assign T_806 = {T_804_1,T_804_0};
  assign T_807 = {T_804_3,T_804_2};
  assign T_808 = {T_807,T_806};
  assign T_809 = {T_804_5,T_804_4};
  assign T_810 = {T_804_7,T_804_6};
  assign T_811 = {T_810,T_809};
  assign T_812 = {T_811,T_808};
  assign T_813 = ~ T_812;
  assign T_814 = timecmp_0 & T_813;
  assign T_815 = T_740 | T_814;
  assign GEN_3 = T_688 ? T_815 : timecmp_0;
  assign GEN_22 = T_661 ? GEN_3 : timecmp_0;
  assign GEN_23 = T_661 ? timecmp_0 : GEN_2;
  assign T_827 = T_658 == 1'h0;
  assign T_828 = T_660 & T_827;
  assign T_848_0 = T_675;
  assign T_860 = T_670 ? T_848_0 : T_692;
  assign T_861 = T_860[0];
  assign T_862 = T_860[1];
  assign T_863 = T_860[2];
  assign T_864 = T_860[3];
  assign T_865 = T_860[4];
  assign T_866 = T_860[5];
  assign T_867 = T_860[6];
  assign T_868 = T_860[7];
  assign GEN_67 = {{7'd0}, T_861};
  assign T_870 = 8'h0 - GEN_67;
  assign T_871 = T_870[7:0];
  assign GEN_68 = {{7'd0}, T_862};
  assign T_873 = 8'h0 - GEN_68;
  assign T_874 = T_873[7:0];
  assign GEN_69 = {{7'd0}, T_863};
  assign T_876 = 8'h0 - GEN_69;
  assign T_877 = T_876[7:0];
  assign GEN_70 = {{7'd0}, T_864};
  assign T_879 = 8'h0 - GEN_70;
  assign T_880 = T_879[7:0];
  assign GEN_71 = {{7'd0}, T_865};
  assign T_882 = 8'h0 - GEN_71;
  assign T_883 = T_882[7:0];
  assign GEN_72 = {{7'd0}, T_866};
  assign T_885 = 8'h0 - GEN_72;
  assign T_886 = T_885[7:0];
  assign GEN_73 = {{7'd0}, T_867};
  assign T_888 = 8'h0 - GEN_73;
  assign T_889 = T_888[7:0];
  assign GEN_74 = {{7'd0}, T_868};
  assign T_891 = 8'h0 - GEN_74;
  assign T_892 = T_891[7:0];
  assign T_898_0 = T_871;
  assign T_898_1 = T_874;
  assign T_898_2 = T_877;
  assign T_898_3 = T_880;
  assign T_898_4 = T_883;
  assign T_898_5 = T_886;
  assign T_898_6 = T_889;
  assign T_898_7 = T_892;
  assign T_900 = {T_898_1,T_898_0};
  assign T_901 = {T_898_3,T_898_2};
  assign T_902 = {T_901,T_900};
  assign T_903 = {T_898_5,T_898_4};
  assign T_904 = {T_898_7,T_898_6};
  assign T_905 = {T_904,T_903};
  assign T_906 = {T_905,T_902};
  assign T_907 = acq_io_deq_bits_data & T_906;
  assign T_921_0 = T_675;
  assign T_933 = T_670 ? T_921_0 : T_692;
  assign T_934 = T_933[0];
  assign T_935 = T_933[1];
  assign T_936 = T_933[2];
  assign T_937 = T_933[3];
  assign T_938 = T_933[4];
  assign T_939 = T_933[5];
  assign T_940 = T_933[6];
  assign T_941 = T_933[7];
  assign GEN_76 = {{7'd0}, T_934};
  assign T_943 = 8'h0 - GEN_76;
  assign T_944 = T_943[7:0];
  assign GEN_77 = {{7'd0}, T_935};
  assign T_946 = 8'h0 - GEN_77;
  assign T_947 = T_946[7:0];
  assign GEN_78 = {{7'd0}, T_936};
  assign T_949 = 8'h0 - GEN_78;
  assign T_950 = T_949[7:0];
  assign GEN_79 = {{7'd0}, T_937};
  assign T_952 = 8'h0 - GEN_79;
  assign T_953 = T_952[7:0];
  assign GEN_80 = {{7'd0}, T_938};
  assign T_955 = 8'h0 - GEN_80;
  assign T_956 = T_955[7:0];
  assign GEN_81 = {{7'd0}, T_939};
  assign T_958 = 8'h0 - GEN_81;
  assign T_959 = T_958[7:0];
  assign GEN_82 = {{7'd0}, T_940};
  assign T_961 = 8'h0 - GEN_82;
  assign T_962 = T_961[7:0];
  assign GEN_83 = {{7'd0}, T_941};
  assign T_964 = 8'h0 - GEN_83;
  assign T_965 = T_964[7:0];
  assign T_971_0 = T_944;
  assign T_971_1 = T_947;
  assign T_971_2 = T_950;
  assign T_971_3 = T_953;
  assign T_971_4 = T_956;
  assign T_971_5 = T_959;
  assign T_971_6 = T_962;
  assign T_971_7 = T_965;
  assign T_973 = {T_971_1,T_971_0};
  assign T_974 = {T_971_3,T_971_2};
  assign T_975 = {T_974,T_973};
  assign T_976 = {T_971_5,T_971_4};
  assign T_977 = {T_971_7,T_971_6};
  assign T_978 = {T_977,T_976};
  assign T_979 = {T_978,T_975};
  assign T_980 = ~ T_979;
  assign GEN_84 = {{32'd0}, ipi_0};
  assign T_981 = GEN_84 & T_980;
  assign T_982 = T_907 | T_981;
  assign GEN_24 = T_688 ? T_982 : {{32'd0}, ipi_0};
  assign T_993 = GEN_84 & 64'h100000001;
  assign GEN_43 = T_828 ? GEN_24 : {{32'd0}, ipi_0};
  assign GEN_44 = T_828 ? T_993 : GEN_23;
  assign T_994 = ipi_0[0];
  assign T_995 = time$ >= timecmp_0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_4 = {2{$random}};
  timecmp_0 = GEN_4[63:0];
  GEN_5 = {2{$random}};
  time$ = GEN_5[63:0];
  GEN_6 = {1{$random}};
  ipi_0 = GEN_6[31:0];
  GEN_7 = {1{$random}};
  GEN_1 = GEN_7[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_661) begin
        if(T_688) begin
          timecmp_0 <= T_815;
        end
      end
    end
    if(reset) begin
      time$ <= 64'h0;
    end else begin
      if(io_rtcTick) begin
        time$ <= T_526;
      end
    end
    if(reset) begin
      ipi_0 <= T_533_0;
    end else begin
      ipi_0 <= GEN_43[31:0];
    end
  end
endmodule
module ROMSlave(
  input   clk,
  input   reset,
  output  io_acquire_ready,
  input   io_acquire_valid,
  input  [25:0] io_acquire_bits_addr_block,
  input  [1:0] io_acquire_bits_client_xact_id,
  input  [2:0] io_acquire_bits_addr_beat,
  input   io_acquire_bits_is_builtin_type,
  input  [2:0] io_acquire_bits_a_type,
  input  [11:0] io_acquire_bits_union,
  input  [63:0] io_acquire_bits_data,
  input   io_grant_ready,
  output  io_grant_valid,
  output [2:0] io_grant_bits_addr_beat,
  output [1:0] io_grant_bits_client_xact_id,
  output  io_grant_bits_manager_xact_id,
  output  io_grant_bits_is_builtin_type,
  output [3:0] io_grant_bits_g_type,
  output [63:0] io_grant_bits_data
);
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_446;
  wire  single_beat;
  wire  T_448;
  wire  multi_beat;
  wire  T_450;
  wire  T_451;
  wire  T_452;
  wire  T_453;
  wire  T_455;
  reg [2:0] addr_beat;
  reg [31:0] GEN_159;
  wire  T_457;
  wire [2:0] GEN_95;
  wire [3:0] T_459;
  wire [2:0] T_460;
  wire [2:0] GEN_1;
  wire  T_461;
  wire [2:0] GEN_2;
  wire [63:0] rom_0;
  wire [63:0] rom_1;
  wire [63:0] rom_2;
  wire [63:0] rom_3;
  wire [63:0] rom_4;
  wire [63:0] rom_5;
  wire [63:0] rom_6;
  wire [63:0] rom_7;
  wire [63:0] rom_8;
  wire [63:0] rom_9;
  wire [63:0] rom_10;
  wire [63:0] rom_11;
  wire [63:0] rom_12;
  wire [63:0] rom_13;
  wire [63:0] rom_14;
  wire [63:0] rom_15;
  wire [63:0] rom_16;
  wire [63:0] rom_17;
  wire [63:0] rom_18;
  wire [63:0] rom_19;
  wire [63:0] rom_20;
  wire [63:0] rom_21;
  wire [63:0] rom_22;
  wire [63:0] rom_23;
  wire [63:0] rom_24;
  wire [63:0] rom_25;
  wire [63:0] rom_26;
  wire [63:0] rom_27;
  wire [63:0] rom_28;
  wire [63:0] rom_29;
  wire [63:0] rom_30;
  wire [63:0] rom_31;
  wire [63:0] rom_32;
  wire [63:0] rom_33;
  wire [63:0] rom_34;
  wire [63:0] rom_35;
  wire [63:0] rom_36;
  wire [63:0] rom_37;
  wire [63:0] rom_38;
  wire [63:0] rom_39;
  wire [63:0] rom_40;
  wire [63:0] rom_41;
  wire [63:0] rom_42;
  wire [63:0] rom_43;
  wire [63:0] rom_44;
  wire [63:0] rom_45;
  wire [63:0] rom_46;
  wire [63:0] rom_47;
  wire [63:0] rom_48;
  wire [63:0] rom_49;
  wire [63:0] rom_50;
  wire [63:0] rom_51;
  wire [63:0] rom_52;
  wire [63:0] rom_53;
  wire [63:0] rom_54;
  wire [63:0] rom_55;
  wire [63:0] rom_56;
  wire [63:0] rom_57;
  wire [63:0] rom_58;
  wire [63:0] rom_59;
  wire [63:0] rom_60;
  wire [63:0] rom_61;
  wire [63:0] rom_62;
  wire [63:0] rom_63;
  wire [63:0] rom_64;
  wire [63:0] rom_65;
  wire [63:0] rom_66;
  wire [63:0] rom_67;
  wire [63:0] rom_68;
  wire [63:0] rom_69;
  wire [63:0] rom_70;
  wire [63:0] rom_71;
  wire [63:0] rom_72;
  wire [63:0] rom_73;
  wire [63:0] rom_74;
  wire [63:0] rom_75;
  wire [63:0] rom_76;
  wire [63:0] rom_77;
  wire [63:0] rom_78;
  wire [63:0] rom_79;
  wire [63:0] rom_80;
  wire [63:0] rom_81;
  wire [63:0] rom_82;
  wire [63:0] rom_83;
  wire [63:0] rom_84;
  wire [63:0] rom_85;
  wire [63:0] rom_86;
  wire [63:0] rom_87;
  wire [63:0] rom_88;
  wire [63:0] rom_89;
  wire [63:0] rom_90;
  wire [63:0] rom_91;
  wire [63:0] rom_92;
  wire [28:0] raddr;
  wire [6:0] T_561;
  wire  T_563;
  wire  T_565;
  wire  last;
  wire  T_566;
  wire  T_583;
  wire [2:0] T_584;
  wire  T_585;
  wire [2:0] T_586;
  wire  T_587;
  wire [2:0] T_588;
  wire  T_589;
  wire [2:0] T_590;
  wire  T_591;
  wire [2:0] T_592;
  wire  T_593;
  wire [2:0] T_594;
  wire  T_595;
  wire [2:0] T_596;
  wire [2:0] T_620_addr_beat;
  wire [1:0] T_620_client_xact_id;
  wire  T_620_manager_xact_id;
  wire  T_620_is_builtin_type;
  wire [3:0] T_620_g_type;
  wire [63:0] T_620_data;
  wire [63:0] GEN_0;
  wire [6:0] GEN_96;
  wire [63:0] GEN_3;
  wire [6:0] GEN_97;
  wire [63:0] GEN_4;
  wire [6:0] GEN_98;
  wire [63:0] GEN_5;
  wire [6:0] GEN_99;
  wire [63:0] GEN_6;
  wire [6:0] GEN_100;
  wire [63:0] GEN_7;
  wire [6:0] GEN_101;
  wire [63:0] GEN_8;
  wire [6:0] GEN_102;
  wire [63:0] GEN_9;
  wire [6:0] GEN_103;
  wire [63:0] GEN_10;
  wire [6:0] GEN_104;
  wire [63:0] GEN_11;
  wire [6:0] GEN_105;
  wire [63:0] GEN_12;
  wire [6:0] GEN_106;
  wire [63:0] GEN_13;
  wire [6:0] GEN_107;
  wire [63:0] GEN_14;
  wire [6:0] GEN_108;
  wire [63:0] GEN_15;
  wire [6:0] GEN_109;
  wire [63:0] GEN_16;
  wire [6:0] GEN_110;
  wire [63:0] GEN_17;
  wire [6:0] GEN_111;
  wire [63:0] GEN_18;
  wire [6:0] GEN_112;
  wire [63:0] GEN_19;
  wire [6:0] GEN_113;
  wire [63:0] GEN_20;
  wire [6:0] GEN_114;
  wire [63:0] GEN_21;
  wire [6:0] GEN_115;
  wire [63:0] GEN_22;
  wire [6:0] GEN_116;
  wire [63:0] GEN_23;
  wire [6:0] GEN_117;
  wire [63:0] GEN_24;
  wire [6:0] GEN_118;
  wire [63:0] GEN_25;
  wire [6:0] GEN_119;
  wire [63:0] GEN_26;
  wire [6:0] GEN_120;
  wire [63:0] GEN_27;
  wire [6:0] GEN_121;
  wire [63:0] GEN_28;
  wire [6:0] GEN_122;
  wire [63:0] GEN_29;
  wire [6:0] GEN_123;
  wire [63:0] GEN_30;
  wire [6:0] GEN_124;
  wire [63:0] GEN_31;
  wire [6:0] GEN_125;
  wire [63:0] GEN_32;
  wire [6:0] GEN_126;
  wire [63:0] GEN_33;
  wire [6:0] GEN_127;
  wire [63:0] GEN_34;
  wire [6:0] GEN_128;
  wire [63:0] GEN_35;
  wire [6:0] GEN_129;
  wire [63:0] GEN_36;
  wire [6:0] GEN_130;
  wire [63:0] GEN_37;
  wire [6:0] GEN_131;
  wire [63:0] GEN_38;
  wire [6:0] GEN_132;
  wire [63:0] GEN_39;
  wire [6:0] GEN_133;
  wire [63:0] GEN_40;
  wire [6:0] GEN_134;
  wire [63:0] GEN_41;
  wire [6:0] GEN_135;
  wire [63:0] GEN_42;
  wire [6:0] GEN_136;
  wire [63:0] GEN_43;
  wire [6:0] GEN_137;
  wire [63:0] GEN_44;
  wire [6:0] GEN_138;
  wire [63:0] GEN_45;
  wire [6:0] GEN_139;
  wire [63:0] GEN_46;
  wire [6:0] GEN_140;
  wire [63:0] GEN_47;
  wire [6:0] GEN_141;
  wire [63:0] GEN_48;
  wire [6:0] GEN_142;
  wire [63:0] GEN_49;
  wire [6:0] GEN_143;
  wire [63:0] GEN_50;
  wire [6:0] GEN_144;
  wire [63:0] GEN_51;
  wire [6:0] GEN_145;
  wire [63:0] GEN_52;
  wire [6:0] GEN_146;
  wire [63:0] GEN_53;
  wire [6:0] GEN_147;
  wire [63:0] GEN_54;
  wire [6:0] GEN_148;
  wire [63:0] GEN_55;
  wire [6:0] GEN_149;
  wire [63:0] GEN_56;
  wire [6:0] GEN_150;
  wire [63:0] GEN_57;
  wire [6:0] GEN_151;
  wire [63:0] GEN_58;
  wire [6:0] GEN_152;
  wire [63:0] GEN_59;
  wire [6:0] GEN_153;
  wire [63:0] GEN_60;
  wire [6:0] GEN_154;
  wire [63:0] GEN_61;
  wire [6:0] GEN_155;
  wire [63:0] GEN_62;
  wire [6:0] GEN_156;
  wire [63:0] GEN_63;
  wire [6:0] GEN_157;
  wire [63:0] GEN_64;
  wire [6:0] GEN_158;
  wire [63:0] GEN_65;
  wire [63:0] GEN_66;
  wire [63:0] GEN_67;
  wire [63:0] GEN_68;
  wire [63:0] GEN_69;
  wire [63:0] GEN_70;
  wire [63:0] GEN_71;
  wire [63:0] GEN_72;
  wire [63:0] GEN_73;
  wire [63:0] GEN_74;
  wire [63:0] GEN_75;
  wire [63:0] GEN_76;
  wire [63:0] GEN_77;
  wire [63:0] GEN_78;
  wire [63:0] GEN_79;
  wire [63:0] GEN_80;
  wire [63:0] GEN_81;
  wire [63:0] GEN_82;
  wire [63:0] GEN_83;
  wire [63:0] GEN_84;
  wire [63:0] GEN_85;
  wire [63:0] GEN_86;
  wire [63:0] GEN_87;
  wire [63:0] GEN_88;
  wire [63:0] GEN_89;
  wire [63:0] GEN_90;
  wire [63:0] GEN_91;
  wire [63:0] GEN_92;
  wire [63:0] GEN_93;
  wire [63:0] GEN_94;
  Queue_20 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_acquire_ready = acq_io_enq_ready;
  assign io_grant_valid = acq_io_deq_valid;
  assign io_grant_bits_addr_beat = T_620_addr_beat;
  assign io_grant_bits_client_xact_id = T_620_client_xact_id;
  assign io_grant_bits_manager_xact_id = T_620_manager_xact_id;
  assign io_grant_bits_is_builtin_type = T_620_is_builtin_type;
  assign io_grant_bits_g_type = T_620_g_type;
  assign io_grant_bits_data = T_620_data;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_acquire_bits_union;
  assign acq_io_enq_bits_data = io_acquire_bits_data;
  assign acq_io_deq_ready = T_566;
  assign T_446 = acq_io_deq_bits_a_type == 3'h0;
  assign single_beat = acq_io_deq_bits_is_builtin_type & T_446;
  assign T_448 = acq_io_deq_bits_a_type == 3'h1;
  assign multi_beat = acq_io_deq_bits_is_builtin_type & T_448;
  assign T_450 = acq_io_deq_valid == 1'h0;
  assign T_451 = T_450 | single_beat;
  assign T_452 = T_451 | multi_beat;
  assign T_453 = T_452 | reset;
  assign T_455 = T_453 == 1'h0;
  assign T_457 = io_grant_ready & io_grant_valid;
  assign GEN_95 = {{2'd0}, 1'h1};
  assign T_459 = addr_beat + GEN_95;
  assign T_460 = T_459[2:0];
  assign GEN_1 = T_457 ? T_460 : addr_beat;
  assign T_461 = io_acquire_ready & io_acquire_valid;
  assign GEN_2 = T_461 ? io_acquire_bits_addr_beat : GEN_1;
  assign rom_0 = 64'hff01011b00004137;
  assign rom_1 = 64'h17370040006f;
  assign rom_2 = 64'h607360306070793;
  assign rom_3 = 64'hc7d7030087a683;
  assign rom_4 = 64'hc7b023000027b7;
  assign rom_5 = 64'he7962300d7a423;
  assign rom_6 = 64'h20604630ff67613;
  assign rom_7 = 64'h6000073700078693;
  assign rom_8 = 64'h87f79300874783;
  assign rom_9 = 64'h168693fe079ce3;
  assign rom_10 = 64'h6c60300c70223;
  assign rom_11 = 64'h6ffe0614e3;
  assign rom_12 = 64'h6f57206f6c6c6548;
  assign rom_13 = 64'ha21646c72;
  assign rom_14 = 64'h0;
  assign rom_15 = 64'h0;
  assign rom_16 = 64'h0;
  assign rom_17 = 64'h0;
  assign rom_18 = 64'h0;
  assign rom_19 = 64'h0;
  assign rom_20 = 64'h0;
  assign rom_21 = 64'h0;
  assign rom_22 = 64'h0;
  assign rom_23 = 64'h0;
  assign rom_24 = 64'h0;
  assign rom_25 = 64'h0;
  assign rom_26 = 64'h0;
  assign rom_27 = 64'h0;
  assign rom_28 = 64'h0;
  assign rom_29 = 64'h0;
  assign rom_30 = 64'h0;
  assign rom_31 = 64'h0;
  assign rom_32 = 64'h200a7b2063696c70;
  assign rom_33 = 64'h7469726f69727020;
  assign rom_34 = 64'h3030303478302079;
  assign rom_35 = 64'h20200a3b30303030;
  assign rom_36 = 64'h20676e69646e6570;
  assign rom_37 = 64'h3031303030347830;
  assign rom_38 = 64'h646e20200a3b3030;
  assign rom_39 = 64'h7d0a3b3220737665;
  assign rom_40 = 64'ha7b206374720a3b;
  assign rom_41 = 64'h3020726464612020;
  assign rom_42 = 64'h6666623030343478;
  assign rom_43 = 64'h61720a3b7d0a3b38;
  assign rom_44 = 64'h203020200a7b206d;
  assign rom_45 = 64'h6461202020200a7b;
  assign rom_46 = 64'h3030387830207264;
  assign rom_47 = 64'h200a3b3030303030;
  assign rom_48 = 64'h20657a6973202020;
  assign rom_49 = 64'h3030303030387830;
  assign rom_50 = 64'h3b7d20200a3b3030;
  assign rom_51 = 64'h65726f630a3b7d0a;
  assign rom_52 = 64'h7b203020200a7b20;
  assign rom_53 = 64'h7b2030202020200a;
  assign rom_54 = 64'h692020202020200a;
  assign rom_55 = 64'h6934367672206173;
  assign rom_56 = 64'h202020200a3b616d;
  assign rom_57 = 64'h6d63656d69742020;
  assign rom_58 = 64'h3030343478302070;
  assign rom_59 = 64'h20200a3b30303034;
  assign rom_60 = 64'h2069706920202020;
  assign rom_61 = 64'h3030303034347830;
  assign rom_62 = 64'h202020200a3b3030;
  assign rom_63 = 64'h7b2063696c702020;
  assign rom_64 = 64'h202020202020200a;
  assign rom_65 = 64'h2020200a7b206d20;
  assign rom_66 = 64'h6569202020202020;
  assign rom_67 = 64'h3230303034783020;
  assign rom_68 = 64'h2020200a3b303030;
  assign rom_69 = 64'h6874202020202020;
  assign rom_70 = 64'h3478302068736572;
  assign rom_71 = 64'h3b30303030303230;
  assign rom_72 = 64'h202020202020200a;
  assign rom_73 = 64'h206d69616c632020;
  assign rom_74 = 64'h3030303230347830;
  assign rom_75 = 64'h202020200a3b3430;
  assign rom_76 = 64'h200a3b7d20202020;
  assign rom_77 = 64'h7320202020202020;
  assign rom_78 = 64'h20202020200a7b20;
  assign rom_79 = 64'h3020656920202020;
  assign rom_80 = 64'h3830323030303478;
  assign rom_81 = 64'h20202020200a3b30;
  assign rom_82 = 64'h6572687420202020;
  assign rom_83 = 64'h3230347830206873;
  assign rom_84 = 64'h200a3b3030303130;
  assign rom_85 = 64'h2020202020202020;
  assign rom_86 = 64'h7830206d69616c63;
  assign rom_87 = 64'h3430303130323034;
  assign rom_88 = 64'h2020202020200a3b;
  assign rom_89 = 64'h2020200a3b7d2020;
  assign rom_90 = 64'h20200a3b7d202020;
  assign rom_91 = 64'h7d20200a3b7d2020;
  assign rom_92 = 64'ha3b7d0a3b;
  assign raddr = {acq_io_deq_bits_addr_block,addr_beat};
  assign T_561 = raddr[6:0];
  assign T_563 = multi_beat == 1'h0;
  assign T_565 = addr_beat == 3'h7;
  assign last = T_563 | T_565;
  assign T_566 = io_grant_ready & last;
  assign T_583 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_584 = T_583 ? 3'h1 : 3'h3;
  assign T_585 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_586 = T_585 ? 3'h1 : T_584;
  assign T_587 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_588 = T_587 ? 3'h4 : T_586;
  assign T_589 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_590 = T_589 ? 3'h3 : T_588;
  assign T_591 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_592 = T_591 ? 3'h3 : T_590;
  assign T_593 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_594 = T_593 ? 3'h5 : T_592;
  assign T_595 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_596 = T_595 ? 3'h4 : T_594;
  assign T_620_addr_beat = addr_beat;
  assign T_620_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_620_manager_xact_id = 1'h0;
  assign T_620_is_builtin_type = 1'h1;
  assign T_620_g_type = {{1'd0}, T_596};
  assign T_620_data = GEN_0;
  assign GEN_0 = GEN_94;
  assign GEN_96 = {{6'd0}, 1'h1};
  assign GEN_3 = GEN_96 == T_561 ? rom_1 : rom_0;
  assign GEN_97 = {{5'd0}, 2'h2};
  assign GEN_4 = GEN_97 == T_561 ? rom_2 : GEN_3;
  assign GEN_98 = {{5'd0}, 2'h3};
  assign GEN_5 = GEN_98 == T_561 ? rom_3 : GEN_4;
  assign GEN_99 = {{4'd0}, 3'h4};
  assign GEN_6 = GEN_99 == T_561 ? rom_4 : GEN_5;
  assign GEN_100 = {{4'd0}, 3'h5};
  assign GEN_7 = GEN_100 == T_561 ? rom_5 : GEN_6;
  assign GEN_101 = {{4'd0}, 3'h6};
  assign GEN_8 = GEN_101 == T_561 ? rom_6 : GEN_7;
  assign GEN_102 = {{4'd0}, 3'h7};
  assign GEN_9 = GEN_102 == T_561 ? rom_7 : GEN_8;
  assign GEN_103 = {{3'd0}, 4'h8};
  assign GEN_10 = GEN_103 == T_561 ? rom_8 : GEN_9;
  assign GEN_104 = {{3'd0}, 4'h9};
  assign GEN_11 = GEN_104 == T_561 ? rom_9 : GEN_10;
  assign GEN_105 = {{3'd0}, 4'ha};
  assign GEN_12 = GEN_105 == T_561 ? rom_10 : GEN_11;
  assign GEN_106 = {{3'd0}, 4'hb};
  assign GEN_13 = GEN_106 == T_561 ? rom_11 : GEN_12;
  assign GEN_107 = {{3'd0}, 4'hc};
  assign GEN_14 = GEN_107 == T_561 ? rom_12 : GEN_13;
  assign GEN_108 = {{3'd0}, 4'hd};
  assign GEN_15 = GEN_108 == T_561 ? rom_13 : GEN_14;
  assign GEN_109 = {{3'd0}, 4'he};
  assign GEN_16 = GEN_109 == T_561 ? rom_14 : GEN_15;
  assign GEN_110 = {{3'd0}, 4'hf};
  assign GEN_17 = GEN_110 == T_561 ? rom_15 : GEN_16;
  assign GEN_111 = {{2'd0}, 5'h10};
  assign GEN_18 = GEN_111 == T_561 ? rom_16 : GEN_17;
  assign GEN_112 = {{2'd0}, 5'h11};
  assign GEN_19 = GEN_112 == T_561 ? rom_17 : GEN_18;
  assign GEN_113 = {{2'd0}, 5'h12};
  assign GEN_20 = GEN_113 == T_561 ? rom_18 : GEN_19;
  assign GEN_114 = {{2'd0}, 5'h13};
  assign GEN_21 = GEN_114 == T_561 ? rom_19 : GEN_20;
  assign GEN_115 = {{2'd0}, 5'h14};
  assign GEN_22 = GEN_115 == T_561 ? rom_20 : GEN_21;
  assign GEN_116 = {{2'd0}, 5'h15};
  assign GEN_23 = GEN_116 == T_561 ? rom_21 : GEN_22;
  assign GEN_117 = {{2'd0}, 5'h16};
  assign GEN_24 = GEN_117 == T_561 ? rom_22 : GEN_23;
  assign GEN_118 = {{2'd0}, 5'h17};
  assign GEN_25 = GEN_118 == T_561 ? rom_23 : GEN_24;
  assign GEN_119 = {{2'd0}, 5'h18};
  assign GEN_26 = GEN_119 == T_561 ? rom_24 : GEN_25;
  assign GEN_120 = {{2'd0}, 5'h19};
  assign GEN_27 = GEN_120 == T_561 ? rom_25 : GEN_26;
  assign GEN_121 = {{2'd0}, 5'h1a};
  assign GEN_28 = GEN_121 == T_561 ? rom_26 : GEN_27;
  assign GEN_122 = {{2'd0}, 5'h1b};
  assign GEN_29 = GEN_122 == T_561 ? rom_27 : GEN_28;
  assign GEN_123 = {{2'd0}, 5'h1c};
  assign GEN_30 = GEN_123 == T_561 ? rom_28 : GEN_29;
  assign GEN_124 = {{2'd0}, 5'h1d};
  assign GEN_31 = GEN_124 == T_561 ? rom_29 : GEN_30;
  assign GEN_125 = {{2'd0}, 5'h1e};
  assign GEN_32 = GEN_125 == T_561 ? rom_30 : GEN_31;
  assign GEN_126 = {{2'd0}, 5'h1f};
  assign GEN_33 = GEN_126 == T_561 ? rom_31 : GEN_32;
  assign GEN_127 = {{1'd0}, 6'h20};
  assign GEN_34 = GEN_127 == T_561 ? rom_32 : GEN_33;
  assign GEN_128 = {{1'd0}, 6'h21};
  assign GEN_35 = GEN_128 == T_561 ? rom_33 : GEN_34;
  assign GEN_129 = {{1'd0}, 6'h22};
  assign GEN_36 = GEN_129 == T_561 ? rom_34 : GEN_35;
  assign GEN_130 = {{1'd0}, 6'h23};
  assign GEN_37 = GEN_130 == T_561 ? rom_35 : GEN_36;
  assign GEN_131 = {{1'd0}, 6'h24};
  assign GEN_38 = GEN_131 == T_561 ? rom_36 : GEN_37;
  assign GEN_132 = {{1'd0}, 6'h25};
  assign GEN_39 = GEN_132 == T_561 ? rom_37 : GEN_38;
  assign GEN_133 = {{1'd0}, 6'h26};
  assign GEN_40 = GEN_133 == T_561 ? rom_38 : GEN_39;
  assign GEN_134 = {{1'd0}, 6'h27};
  assign GEN_41 = GEN_134 == T_561 ? rom_39 : GEN_40;
  assign GEN_135 = {{1'd0}, 6'h28};
  assign GEN_42 = GEN_135 == T_561 ? rom_40 : GEN_41;
  assign GEN_136 = {{1'd0}, 6'h29};
  assign GEN_43 = GEN_136 == T_561 ? rom_41 : GEN_42;
  assign GEN_137 = {{1'd0}, 6'h2a};
  assign GEN_44 = GEN_137 == T_561 ? rom_42 : GEN_43;
  assign GEN_138 = {{1'd0}, 6'h2b};
  assign GEN_45 = GEN_138 == T_561 ? rom_43 : GEN_44;
  assign GEN_139 = {{1'd0}, 6'h2c};
  assign GEN_46 = GEN_139 == T_561 ? rom_44 : GEN_45;
  assign GEN_140 = {{1'd0}, 6'h2d};
  assign GEN_47 = GEN_140 == T_561 ? rom_45 : GEN_46;
  assign GEN_141 = {{1'd0}, 6'h2e};
  assign GEN_48 = GEN_141 == T_561 ? rom_46 : GEN_47;
  assign GEN_142 = {{1'd0}, 6'h2f};
  assign GEN_49 = GEN_142 == T_561 ? rom_47 : GEN_48;
  assign GEN_143 = {{1'd0}, 6'h30};
  assign GEN_50 = GEN_143 == T_561 ? rom_48 : GEN_49;
  assign GEN_144 = {{1'd0}, 6'h31};
  assign GEN_51 = GEN_144 == T_561 ? rom_49 : GEN_50;
  assign GEN_145 = {{1'd0}, 6'h32};
  assign GEN_52 = GEN_145 == T_561 ? rom_50 : GEN_51;
  assign GEN_146 = {{1'd0}, 6'h33};
  assign GEN_53 = GEN_146 == T_561 ? rom_51 : GEN_52;
  assign GEN_147 = {{1'd0}, 6'h34};
  assign GEN_54 = GEN_147 == T_561 ? rom_52 : GEN_53;
  assign GEN_148 = {{1'd0}, 6'h35};
  assign GEN_55 = GEN_148 == T_561 ? rom_53 : GEN_54;
  assign GEN_149 = {{1'd0}, 6'h36};
  assign GEN_56 = GEN_149 == T_561 ? rom_54 : GEN_55;
  assign GEN_150 = {{1'd0}, 6'h37};
  assign GEN_57 = GEN_150 == T_561 ? rom_55 : GEN_56;
  assign GEN_151 = {{1'd0}, 6'h38};
  assign GEN_58 = GEN_151 == T_561 ? rom_56 : GEN_57;
  assign GEN_152 = {{1'd0}, 6'h39};
  assign GEN_59 = GEN_152 == T_561 ? rom_57 : GEN_58;
  assign GEN_153 = {{1'd0}, 6'h3a};
  assign GEN_60 = GEN_153 == T_561 ? rom_58 : GEN_59;
  assign GEN_154 = {{1'd0}, 6'h3b};
  assign GEN_61 = GEN_154 == T_561 ? rom_59 : GEN_60;
  assign GEN_155 = {{1'd0}, 6'h3c};
  assign GEN_62 = GEN_155 == T_561 ? rom_60 : GEN_61;
  assign GEN_156 = {{1'd0}, 6'h3d};
  assign GEN_63 = GEN_156 == T_561 ? rom_61 : GEN_62;
  assign GEN_157 = {{1'd0}, 6'h3e};
  assign GEN_64 = GEN_157 == T_561 ? rom_62 : GEN_63;
  assign GEN_158 = {{1'd0}, 6'h3f};
  assign GEN_65 = GEN_158 == T_561 ? rom_63 : GEN_64;
  assign GEN_66 = 7'h40 == T_561 ? rom_64 : GEN_65;
  assign GEN_67 = 7'h41 == T_561 ? rom_65 : GEN_66;
  assign GEN_68 = 7'h42 == T_561 ? rom_66 : GEN_67;
  assign GEN_69 = 7'h43 == T_561 ? rom_67 : GEN_68;
  assign GEN_70 = 7'h44 == T_561 ? rom_68 : GEN_69;
  assign GEN_71 = 7'h45 == T_561 ? rom_69 : GEN_70;
  assign GEN_72 = 7'h46 == T_561 ? rom_70 : GEN_71;
  assign GEN_73 = 7'h47 == T_561 ? rom_71 : GEN_72;
  assign GEN_74 = 7'h48 == T_561 ? rom_72 : GEN_73;
  assign GEN_75 = 7'h49 == T_561 ? rom_73 : GEN_74;
  assign GEN_76 = 7'h4a == T_561 ? rom_74 : GEN_75;
  assign GEN_77 = 7'h4b == T_561 ? rom_75 : GEN_76;
  assign GEN_78 = 7'h4c == T_561 ? rom_76 : GEN_77;
  assign GEN_79 = 7'h4d == T_561 ? rom_77 : GEN_78;
  assign GEN_80 = 7'h4e == T_561 ? rom_78 : GEN_79;
  assign GEN_81 = 7'h4f == T_561 ? rom_79 : GEN_80;
  assign GEN_82 = 7'h50 == T_561 ? rom_80 : GEN_81;
  assign GEN_83 = 7'h51 == T_561 ? rom_81 : GEN_82;
  assign GEN_84 = 7'h52 == T_561 ? rom_82 : GEN_83;
  assign GEN_85 = 7'h53 == T_561 ? rom_83 : GEN_84;
  assign GEN_86 = 7'h54 == T_561 ? rom_84 : GEN_85;
  assign GEN_87 = 7'h55 == T_561 ? rom_85 : GEN_86;
  assign GEN_88 = 7'h56 == T_561 ? rom_86 : GEN_87;
  assign GEN_89 = 7'h57 == T_561 ? rom_87 : GEN_88;
  assign GEN_90 = 7'h58 == T_561 ? rom_88 : GEN_89;
  assign GEN_91 = 7'h59 == T_561 ? rom_89 : GEN_90;
  assign GEN_92 = 7'h5a == T_561 ? rom_90 : GEN_91;
  assign GEN_93 = 7'h5b == T_561 ? rom_91 : GEN_92;
  assign GEN_94 = 7'h5c == T_561 ? rom_92 : GEN_93;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_159 = {1{$random}};
  addr_beat = GEN_159[2:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_461) begin
        addr_beat <= io_acquire_bits_addr_beat;
      end else begin
        if(T_457) begin
          addr_beat <= T_460;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_455) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported ROMSlave operation\n    at Rom.scala:17 assert(!acq.valid || single_beat || multi_beat, \"unsupported ROMSlave operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_455) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_455) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BRAMSlave(
  input   clk,
  input   reset,
  output  io_acquire_ready,
  input   io_acquire_valid,
  input  [25:0] io_acquire_bits_addr_block,
  input  [1:0] io_acquire_bits_client_xact_id,
  input  [2:0] io_acquire_bits_addr_beat,
  input   io_acquire_bits_is_builtin_type,
  input  [2:0] io_acquire_bits_a_type,
  input  [11:0] io_acquire_bits_union,
  input  [63:0] io_acquire_bits_data,
  input   io_grant_ready,
  output  io_grant_valid,
  output [2:0] io_grant_bits_addr_beat,
  output [1:0] io_grant_bits_client_xact_id,
  output  io_grant_bits_manager_xact_id,
  output  io_grant_bits_is_builtin_type,
  output [3:0] io_grant_bits_g_type,
  output [63:0] io_grant_bits_data
);
  reg [7:0] bram_0 [0:8191];
  reg [31:0] GEN_21;
  wire [7:0] bram_0_rdata_data;
  wire [12:0] bram_0_rdata_addr;
  wire  bram_0_rdata_en;
  reg [12:0] GEN_22;
  reg [31:0] GEN_23;
  reg  GEN_24;
  reg [31:0] GEN_25;
  wire [7:0] bram_0_T_767_data;
  wire [12:0] bram_0_T_767_addr;
  wire  bram_0_T_767_mask;
  wire  bram_0_T_767_en;
  reg [7:0] bram_1 [0:8191];
  reg [31:0] GEN_26;
  wire [7:0] bram_1_rdata_data;
  wire [12:0] bram_1_rdata_addr;
  wire  bram_1_rdata_en;
  reg [12:0] GEN_27;
  reg [31:0] GEN_28;
  reg  GEN_29;
  reg [31:0] GEN_30;
  wire [7:0] bram_1_T_767_data;
  wire [12:0] bram_1_T_767_addr;
  wire  bram_1_T_767_mask;
  wire  bram_1_T_767_en;
  reg [7:0] bram_2 [0:8191];
  reg [31:0] GEN_31;
  wire [7:0] bram_2_rdata_data;
  wire [12:0] bram_2_rdata_addr;
  wire  bram_2_rdata_en;
  reg [12:0] GEN_32;
  reg [31:0] GEN_33;
  reg  GEN_34;
  reg [31:0] GEN_35;
  wire [7:0] bram_2_T_767_data;
  wire [12:0] bram_2_T_767_addr;
  wire  bram_2_T_767_mask;
  wire  bram_2_T_767_en;
  reg [7:0] bram_3 [0:8191];
  reg [31:0] GEN_36;
  wire [7:0] bram_3_rdata_data;
  wire [12:0] bram_3_rdata_addr;
  wire  bram_3_rdata_en;
  reg [12:0] GEN_37;
  reg [31:0] GEN_38;
  reg  GEN_39;
  reg [31:0] GEN_40;
  wire [7:0] bram_3_T_767_data;
  wire [12:0] bram_3_T_767_addr;
  wire  bram_3_T_767_mask;
  wire  bram_3_T_767_en;
  reg [7:0] bram_4 [0:8191];
  reg [31:0] GEN_41;
  wire [7:0] bram_4_rdata_data;
  wire [12:0] bram_4_rdata_addr;
  wire  bram_4_rdata_en;
  reg [12:0] GEN_43;
  reg [31:0] GEN_45;
  reg  GEN_47;
  reg [31:0] GEN_49;
  wire [7:0] bram_4_T_767_data;
  wire [12:0] bram_4_T_767_addr;
  wire  bram_4_T_767_mask;
  wire  bram_4_T_767_en;
  reg [7:0] bram_5 [0:8191];
  reg [31:0] GEN_51;
  wire [7:0] bram_5_rdata_data;
  wire [12:0] bram_5_rdata_addr;
  wire  bram_5_rdata_en;
  reg [12:0] GEN_53;
  reg [31:0] GEN_55;
  reg  GEN_58;
  reg [31:0] GEN_60;
  wire [7:0] bram_5_T_767_data;
  wire [12:0] bram_5_T_767_addr;
  wire  bram_5_T_767_mask;
  wire  bram_5_T_767_en;
  reg [7:0] bram_6 [0:8191];
  reg [31:0] GEN_61;
  wire [7:0] bram_6_rdata_data;
  wire [12:0] bram_6_rdata_addr;
  wire  bram_6_rdata_en;
  reg [12:0] GEN_64;
  reg [31:0] GEN_65;
  reg  GEN_66;
  reg [31:0] GEN_67;
  wire [7:0] bram_6_T_767_data;
  wire [12:0] bram_6_T_767_addr;
  wire  bram_6_T_767_mask;
  wire  bram_6_T_767_en;
  reg [7:0] bram_7 [0:8191];
  reg [31:0] GEN_68;
  wire [7:0] bram_7_rdata_data;
  wire [12:0] bram_7_rdata_addr;
  wire  bram_7_rdata_en;
  reg [12:0] GEN_69;
  reg [31:0] GEN_70;
  reg  GEN_71;
  reg [31:0] GEN_72;
  wire [7:0] bram_7_T_767_data;
  wire [12:0] bram_7_T_767_addr;
  wire  bram_7_T_767_mask;
  wire  bram_7_T_767_en;
  reg [1:0] state;
  reg [31:0] GEN_73;
  reg [25:0] r_acq_addr_block;
  reg [31:0] GEN_74;
  reg [1:0] r_acq_client_xact_id;
  reg [31:0] GEN_75;
  reg [2:0] r_acq_addr_beat;
  reg [31:0] GEN_76;
  reg  r_acq_is_builtin_type;
  reg [31:0] GEN_77;
  reg [2:0] r_acq_a_type;
  reg [31:0] GEN_78;
  reg [11:0] r_acq_union;
  reg [31:0] GEN_79;
  wire  T_477;
  wire  is_get;
  wire  T_478;
  wire  is_getblk;
  wire  T_479;
  wire  is_put;
  wire  T_480;
  wire  is_putblk;
  reg [2:0] beats;
  reg [31:0] GEN_80;
  wire  T_482;
  wire  T_483;
  wire  T_485;
  wire  T_487;
  wire  T_488;
  wire  T_489;
  wire  T_490;
  wire [1:0] GEN_0;
  wire [2:0] GEN_1;
  wire [1:0] GEN_2;
  wire [2:0] GEN_3;
  wire [1:0] GEN_4;
  wire [25:0] GEN_5;
  wire [1:0] GEN_6;
  wire [2:0] GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [11:0] GEN_10;
  wire [1:0] GEN_11;
  wire [2:0] GEN_12;
  wire  T_493;
  wire  T_494;
  wire [2:0] GEN_57;
  wire [3:0] T_496;
  wire [2:0] T_497;
  wire [3:0] T_499;
  wire [2:0] T_500;
  wire [2:0] GEN_59;
  wire  T_502;
  wire [1:0] GEN_13;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire [1:0] GEN_16;
  wire  T_503;
  wire  T_504;
  wire [1:0] GEN_17;
  wire [2:0] GEN_18;
  wire [1:0] GEN_19;
  wire  T_510;
  wire  T_511;
  wire [1:0] GEN_20;
  wire [28:0] acq_addr;
  wire [28:0] r_acq_addr;
  wire  T_517;
  wire [28:0] GEN_62;
  wire [29:0] T_519;
  wire [28:0] T_520;
  wire [28:0] T_521;
  wire [28:0] raddr;
  wire [28:0] T_523;
  wire  T_528;
  wire  wen;
  wire [7:0] T_529;
  wire [7:0] T_530;
  wire [7:0] T_531;
  wire [7:0] T_532;
  wire [7:0] T_533;
  wire [7:0] T_534;
  wire [7:0] T_535;
  wire [7:0] T_536;
  wire [7:0] wdata_0;
  wire [7:0] wdata_1;
  wire [7:0] wdata_2;
  wire [7:0] wdata_3;
  wire [7:0] wdata_4;
  wire [7:0] wdata_5;
  wire [7:0] wdata_6;
  wire [7:0] wdata_7;
  wire  T_544;
  wire  T_545;
  wire [7:0] GEN_63;
  wire [8:0] T_549;
  wire [7:0] T_550;
  wire [7:0] T_556_0;
  wire  T_564;
  wire [7:0] T_565;
  wire [7:0] T_567;
  wire [7:0] T_568;
  wire  T_569;
  wire [7:0] T_583_0;
  wire [7:0] T_595;
  wire  T_596;
  wire [7:0] T_610_0;
  wire [7:0] T_622;
  wire  T_623;
  wire [7:0] T_637_0;
  wire [7:0] T_649;
  wire  T_650;
  wire [7:0] T_664_0;
  wire [7:0] T_676;
  wire  T_677;
  wire [7:0] T_691_0;
  wire [7:0] T_703;
  wire  T_704;
  wire [7:0] T_718_0;
  wire [7:0] T_730;
  wire  T_731;
  wire [7:0] T_745_0;
  wire [7:0] T_757;
  wire  T_758;
  wire  wmask_0;
  wire  wmask_1;
  wire  wmask_2;
  wire  wmask_3;
  wire  wmask_4;
  wire  wmask_5;
  wire  wmask_6;
  wire  wmask_7;
  wire  GEN_42;
  wire  GEN_44;
  wire  GEN_46;
  wire  GEN_48;
  wire  GEN_50;
  wire  GEN_52;
  wire  GEN_54;
  wire  GEN_56;
  wire  T_771;
  wire  T_788;
  wire [2:0] T_789;
  wire  T_790;
  wire [2:0] T_791;
  wire  T_792;
  wire [2:0] T_793;
  wire  T_794;
  wire [2:0] T_795;
  wire  T_796;
  wire [2:0] T_797;
  wire  T_798;
  wire [2:0] T_799;
  wire  T_800;
  wire [2:0] T_801;
  wire [15:0] T_803;
  wire [15:0] T_804;
  wire [31:0] T_805;
  wire [15:0] T_806;
  wire [15:0] T_807;
  wire [31:0] T_808;
  wire [63:0] T_809;
  wire [2:0] T_832_addr_beat;
  wire [1:0] T_832_client_xact_id;
  wire  T_832_manager_xact_id;
  wire  T_832_is_builtin_type;
  wire [3:0] T_832_g_type;
  wire [63:0] T_832_data;
  wire  T_856;
  assign io_acquire_ready = T_856;
  assign io_grant_valid = T_771;
  assign io_grant_bits_addr_beat = T_832_addr_beat;
  assign io_grant_bits_client_xact_id = T_832_client_xact_id;
  assign io_grant_bits_manager_xact_id = T_832_manager_xact_id;
  assign io_grant_bits_is_builtin_type = T_832_is_builtin_type;
  assign io_grant_bits_g_type = T_832_g_type;
  assign io_grant_bits_data = T_832_data;
  assign bram_0_rdata_addr = T_523[12:0];
  assign bram_0_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign bram_0_rdata_data = bram_0[GEN_22];
  `else
  assign bram_0_rdata_data = GEN_22 >= 14'h2000 ? $random : bram_0[GEN_22];
  `endif
  assign bram_0_T_767_data = wdata_0;
  assign bram_0_T_767_addr = acq_addr[12:0];
  assign bram_0_T_767_mask = GEN_42;
  assign bram_0_T_767_en = wen;
  assign bram_1_rdata_addr = T_523[12:0];
  assign bram_1_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign bram_1_rdata_data = bram_1[GEN_27];
  `else
  assign bram_1_rdata_data = GEN_27 >= 14'h2000 ? $random : bram_1[GEN_27];
  `endif
  assign bram_1_T_767_data = wdata_1;
  assign bram_1_T_767_addr = acq_addr[12:0];
  assign bram_1_T_767_mask = GEN_44;
  assign bram_1_T_767_en = wen;
  assign bram_2_rdata_addr = T_523[12:0];
  assign bram_2_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign bram_2_rdata_data = bram_2[GEN_32];
  `else
  assign bram_2_rdata_data = GEN_32 >= 14'h2000 ? $random : bram_2[GEN_32];
  `endif
  assign bram_2_T_767_data = wdata_2;
  assign bram_2_T_767_addr = acq_addr[12:0];
  assign bram_2_T_767_mask = GEN_46;
  assign bram_2_T_767_en = wen;
  assign bram_3_rdata_addr = T_523[12:0];
  assign bram_3_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign bram_3_rdata_data = bram_3[GEN_37];
  `else
  assign bram_3_rdata_data = GEN_37 >= 14'h2000 ? $random : bram_3[GEN_37];
  `endif
  assign bram_3_T_767_data = wdata_3;
  assign bram_3_T_767_addr = acq_addr[12:0];
  assign bram_3_T_767_mask = GEN_48;
  assign bram_3_T_767_en = wen;
  assign bram_4_rdata_addr = T_523[12:0];
  assign bram_4_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign bram_4_rdata_data = bram_4[GEN_43];
  `else
  assign bram_4_rdata_data = GEN_43 >= 14'h2000 ? $random : bram_4[GEN_43];
  `endif
  assign bram_4_T_767_data = wdata_4;
  assign bram_4_T_767_addr = acq_addr[12:0];
  assign bram_4_T_767_mask = GEN_50;
  assign bram_4_T_767_en = wen;
  assign bram_5_rdata_addr = T_523[12:0];
  assign bram_5_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign bram_5_rdata_data = bram_5[GEN_53];
  `else
  assign bram_5_rdata_data = GEN_53 >= 14'h2000 ? $random : bram_5[GEN_53];
  `endif
  assign bram_5_T_767_data = wdata_5;
  assign bram_5_T_767_addr = acq_addr[12:0];
  assign bram_5_T_767_mask = GEN_52;
  assign bram_5_T_767_en = wen;
  assign bram_6_rdata_addr = T_523[12:0];
  assign bram_6_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign bram_6_rdata_data = bram_6[GEN_64];
  `else
  assign bram_6_rdata_data = GEN_64 >= 14'h2000 ? $random : bram_6[GEN_64];
  `endif
  assign bram_6_T_767_data = wdata_6;
  assign bram_6_T_767_addr = acq_addr[12:0];
  assign bram_6_T_767_mask = GEN_54;
  assign bram_6_T_767_en = wen;
  assign bram_7_rdata_addr = T_523[12:0];
  assign bram_7_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign bram_7_rdata_data = bram_7[GEN_69];
  `else
  assign bram_7_rdata_data = GEN_69 >= 14'h2000 ? $random : bram_7[GEN_69];
  `endif
  assign bram_7_T_767_data = wdata_7;
  assign bram_7_T_767_addr = acq_addr[12:0];
  assign bram_7_T_767_mask = GEN_56;
  assign bram_7_T_767_en = wen;
  assign T_477 = io_acquire_bits_a_type == 3'h0;
  assign is_get = io_acquire_bits_is_builtin_type & T_477;
  assign T_478 = io_acquire_bits_a_type == 3'h1;
  assign is_getblk = io_acquire_bits_is_builtin_type & T_478;
  assign T_479 = io_acquire_bits_a_type == 3'h2;
  assign is_put = io_acquire_bits_is_builtin_type & T_479;
  assign T_480 = io_acquire_bits_a_type == 3'h3;
  assign is_putblk = io_acquire_bits_is_builtin_type & T_480;
  assign T_482 = io_acquire_ready & io_acquire_valid;
  assign T_483 = is_get | is_put;
  assign T_485 = io_acquire_bits_a_type == 3'h5;
  assign T_487 = io_acquire_bits_a_type == 3'h6;
  assign T_488 = T_485 | T_487;
  assign T_489 = io_acquire_bits_is_builtin_type & T_488;
  assign T_490 = T_483 | T_489;
  assign GEN_0 = T_490 ? 2'h3 : state;
  assign GEN_1 = is_getblk ? 3'h7 : beats;
  assign GEN_2 = is_getblk ? 2'h1 : GEN_0;
  assign GEN_3 = is_putblk ? 3'h6 : GEN_1;
  assign GEN_4 = is_putblk ? 2'h2 : GEN_2;
  assign GEN_5 = T_482 ? io_acquire_bits_addr_block : r_acq_addr_block;
  assign GEN_6 = T_482 ? io_acquire_bits_client_xact_id : r_acq_client_xact_id;
  assign GEN_7 = T_482 ? io_acquire_bits_addr_beat : r_acq_addr_beat;
  assign GEN_8 = T_482 ? io_acquire_bits_is_builtin_type : r_acq_is_builtin_type;
  assign GEN_9 = T_482 ? io_acquire_bits_a_type : r_acq_a_type;
  assign GEN_10 = T_482 ? io_acquire_bits_union : r_acq_union;
  assign GEN_11 = T_482 ? GEN_4 : state;
  assign GEN_12 = T_482 ? GEN_3 : beats;
  assign T_493 = state == 2'h1;
  assign T_494 = T_493 & io_grant_ready;
  assign GEN_57 = {{2'd0}, 1'h1};
  assign T_496 = r_acq_addr_beat + GEN_57;
  assign T_497 = T_496[2:0];
  assign T_499 = beats - GEN_57;
  assign T_500 = T_499[2:0];
  assign GEN_59 = {{2'd0}, 1'h0};
  assign T_502 = beats == GEN_59;
  assign GEN_13 = T_502 ? 2'h0 : GEN_11;
  assign GEN_14 = T_494 ? T_497 : GEN_7;
  assign GEN_15 = T_494 ? T_500 : GEN_12;
  assign GEN_16 = T_494 ? GEN_13 : GEN_11;
  assign T_503 = state == 2'h2;
  assign T_504 = T_503 & io_acquire_valid;
  assign GEN_17 = T_502 ? 2'h3 : GEN_16;
  assign GEN_18 = T_504 ? T_500 : GEN_15;
  assign GEN_19 = T_504 ? GEN_17 : GEN_16;
  assign T_510 = state == 2'h3;
  assign T_511 = T_510 & io_grant_ready;
  assign GEN_20 = T_511 ? 2'h0 : GEN_19;
  assign acq_addr = {io_acquire_bits_addr_block,io_acquire_bits_addr_beat};
  assign r_acq_addr = {r_acq_addr_block,r_acq_addr_beat};
  assign T_517 = state == 2'h0;
  assign GEN_62 = {{28'd0}, 1'h1};
  assign T_519 = r_acq_addr + GEN_62;
  assign T_520 = T_519[28:0];
  assign T_521 = io_grant_ready ? T_520 : r_acq_addr;
  assign raddr = T_517 ? acq_addr : T_521;
  assign T_523 = raddr;
  assign T_528 = is_put | is_putblk;
  assign wen = T_482 & T_528;
  assign T_529 = io_acquire_bits_data[7:0];
  assign T_530 = io_acquire_bits_data[15:8];
  assign T_531 = io_acquire_bits_data[23:16];
  assign T_532 = io_acquire_bits_data[31:24];
  assign T_533 = io_acquire_bits_data[39:32];
  assign T_534 = io_acquire_bits_data[47:40];
  assign T_535 = io_acquire_bits_data[55:48];
  assign T_536 = io_acquire_bits_data[63:56];
  assign wdata_0 = T_529;
  assign wdata_1 = T_530;
  assign wdata_2 = T_531;
  assign wdata_3 = T_532;
  assign wdata_4 = T_533;
  assign wdata_5 = T_534;
  assign wdata_6 = T_535;
  assign wdata_7 = T_536;
  assign T_544 = io_acquire_bits_a_type == 3'h4;
  assign T_545 = io_acquire_bits_is_builtin_type & T_544;
  assign GEN_63 = {{7'd0}, 1'h1};
  assign T_549 = 8'h0 - GEN_63;
  assign T_550 = T_549[7:0];
  assign T_556_0 = T_550;
  assign T_564 = is_putblk | is_put;
  assign T_565 = io_acquire_bits_union[8:1];
  assign T_567 = T_564 ? T_565 : {{7'd0}, 1'h0};
  assign T_568 = T_545 ? T_556_0 : T_567;
  assign T_569 = T_568[0];
  assign T_583_0 = T_550;
  assign T_595 = T_545 ? T_583_0 : T_567;
  assign T_596 = T_595[1];
  assign T_610_0 = T_550;
  assign T_622 = T_545 ? T_610_0 : T_567;
  assign T_623 = T_622[2];
  assign T_637_0 = T_550;
  assign T_649 = T_545 ? T_637_0 : T_567;
  assign T_650 = T_649[3];
  assign T_664_0 = T_550;
  assign T_676 = T_545 ? T_664_0 : T_567;
  assign T_677 = T_676[4];
  assign T_691_0 = T_550;
  assign T_703 = T_545 ? T_691_0 : T_567;
  assign T_704 = T_703[5];
  assign T_718_0 = T_550;
  assign T_730 = T_545 ? T_718_0 : T_567;
  assign T_731 = T_730[6];
  assign T_745_0 = T_550;
  assign T_757 = T_545 ? T_745_0 : T_567;
  assign T_758 = T_757[7];
  assign wmask_0 = T_569;
  assign wmask_1 = T_596;
  assign wmask_2 = T_623;
  assign wmask_3 = T_650;
  assign wmask_4 = T_677;
  assign wmask_5 = T_704;
  assign wmask_6 = T_731;
  assign wmask_7 = T_758;
  assign GEN_42 = wen ? wmask_0 : 1'h0;
  assign GEN_44 = wen ? wmask_1 : 1'h0;
  assign GEN_46 = wen ? wmask_2 : 1'h0;
  assign GEN_48 = wen ? wmask_3 : 1'h0;
  assign GEN_50 = wen ? wmask_4 : 1'h0;
  assign GEN_52 = wen ? wmask_5 : 1'h0;
  assign GEN_54 = wen ? wmask_6 : 1'h0;
  assign GEN_56 = wen ? wmask_7 : 1'h0;
  assign T_771 = T_510 | T_493;
  assign T_788 = 3'h6 == r_acq_a_type;
  assign T_789 = T_788 ? 3'h1 : 3'h3;
  assign T_790 = 3'h5 == r_acq_a_type;
  assign T_791 = T_790 ? 3'h1 : T_789;
  assign T_792 = 3'h4 == r_acq_a_type;
  assign T_793 = T_792 ? 3'h4 : T_791;
  assign T_794 = 3'h3 == r_acq_a_type;
  assign T_795 = T_794 ? 3'h3 : T_793;
  assign T_796 = 3'h2 == r_acq_a_type;
  assign T_797 = T_796 ? 3'h3 : T_795;
  assign T_798 = 3'h1 == r_acq_a_type;
  assign T_799 = T_798 ? 3'h5 : T_797;
  assign T_800 = 3'h0 == r_acq_a_type;
  assign T_801 = T_800 ? 3'h4 : T_799;
  assign T_803 = {bram_1_rdata_data,bram_0_rdata_data};
  assign T_804 = {bram_3_rdata_data,bram_2_rdata_data};
  assign T_805 = {T_804,T_803};
  assign T_806 = {bram_5_rdata_data,bram_4_rdata_data};
  assign T_807 = {bram_7_rdata_data,bram_6_rdata_data};
  assign T_808 = {T_807,T_806};
  assign T_809 = {T_808,T_805};
  assign T_832_addr_beat = r_acq_addr_beat;
  assign T_832_client_xact_id = r_acq_client_xact_id;
  assign T_832_manager_xact_id = 1'h0;
  assign T_832_is_builtin_type = 1'h1;
  assign T_832_g_type = {{1'd0}, T_801};
  assign T_832_data = T_809;
  assign T_856 = T_517 | T_503;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_21 = {1{$random}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    bram_0[initvar] = GEN_21[7:0];
  GEN_23 = {1{$random}};
  GEN_22 = GEN_23[12:0];
  GEN_25 = {1{$random}};
  GEN_24 = GEN_25[0:0];
  GEN_26 = {1{$random}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    bram_1[initvar] = GEN_26[7:0];
  GEN_28 = {1{$random}};
  GEN_27 = GEN_28[12:0];
  GEN_30 = {1{$random}};
  GEN_29 = GEN_30[0:0];
  GEN_31 = {1{$random}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    bram_2[initvar] = GEN_31[7:0];
  GEN_33 = {1{$random}};
  GEN_32 = GEN_33[12:0];
  GEN_35 = {1{$random}};
  GEN_34 = GEN_35[0:0];
  GEN_36 = {1{$random}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    bram_3[initvar] = GEN_36[7:0];
  GEN_38 = {1{$random}};
  GEN_37 = GEN_38[12:0];
  GEN_40 = {1{$random}};
  GEN_39 = GEN_40[0:0];
  GEN_41 = {1{$random}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    bram_4[initvar] = GEN_41[7:0];
  GEN_45 = {1{$random}};
  GEN_43 = GEN_45[12:0];
  GEN_49 = {1{$random}};
  GEN_47 = GEN_49[0:0];
  GEN_51 = {1{$random}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    bram_5[initvar] = GEN_51[7:0];
  GEN_55 = {1{$random}};
  GEN_53 = GEN_55[12:0];
  GEN_60 = {1{$random}};
  GEN_58 = GEN_60[0:0];
  GEN_61 = {1{$random}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    bram_6[initvar] = GEN_61[7:0];
  GEN_65 = {1{$random}};
  GEN_64 = GEN_65[12:0];
  GEN_67 = {1{$random}};
  GEN_66 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    bram_7[initvar] = GEN_68[7:0];
  GEN_70 = {1{$random}};
  GEN_69 = GEN_70[12:0];
  GEN_72 = {1{$random}};
  GEN_71 = GEN_72[0:0];
  GEN_73 = {1{$random}};
  state = GEN_73[1:0];
  GEN_74 = {1{$random}};
  r_acq_addr_block = GEN_74[25:0];
  GEN_75 = {1{$random}};
  r_acq_client_xact_id = GEN_75[1:0];
  GEN_76 = {1{$random}};
  r_acq_addr_beat = GEN_76[2:0];
  GEN_77 = {1{$random}};
  r_acq_is_builtin_type = GEN_77[0:0];
  GEN_78 = {1{$random}};
  r_acq_a_type = GEN_78[2:0];
  GEN_79 = {1{$random}};
  r_acq_union = GEN_79[11:0];
  GEN_80 = {1{$random}};
  beats = GEN_80[2:0];
  end
`endif
  always @(posedge clk) begin
    GEN_22 <= bram_0_rdata_addr;
    GEN_24 <= bram_0_rdata_en;
    if(bram_0_T_767_en & bram_0_T_767_mask) begin
      bram_0[bram_0_T_767_addr] <= bram_0_T_767_data;
    end
    GEN_27 <= bram_1_rdata_addr;
    GEN_29 <= bram_1_rdata_en;
    if(bram_1_T_767_en & bram_1_T_767_mask) begin
      bram_1[bram_1_T_767_addr] <= bram_1_T_767_data;
    end
    GEN_32 <= bram_2_rdata_addr;
    GEN_34 <= bram_2_rdata_en;
    if(bram_2_T_767_en & bram_2_T_767_mask) begin
      bram_2[bram_2_T_767_addr] <= bram_2_T_767_data;
    end
    GEN_37 <= bram_3_rdata_addr;
    GEN_39 <= bram_3_rdata_en;
    if(bram_3_T_767_en & bram_3_T_767_mask) begin
      bram_3[bram_3_T_767_addr] <= bram_3_T_767_data;
    end
    GEN_43 <= bram_4_rdata_addr;
    GEN_47 <= bram_4_rdata_en;
    if(bram_4_T_767_en & bram_4_T_767_mask) begin
      bram_4[bram_4_T_767_addr] <= bram_4_T_767_data;
    end
    GEN_53 <= bram_5_rdata_addr;
    GEN_58 <= bram_5_rdata_en;
    if(bram_5_T_767_en & bram_5_T_767_mask) begin
      bram_5[bram_5_T_767_addr] <= bram_5_T_767_data;
    end
    GEN_64 <= bram_6_rdata_addr;
    GEN_66 <= bram_6_rdata_en;
    if(bram_6_T_767_en & bram_6_T_767_mask) begin
      bram_6[bram_6_T_767_addr] <= bram_6_T_767_data;
    end
    GEN_69 <= bram_7_rdata_addr;
    GEN_71 <= bram_7_rdata_en;
    if(bram_7_T_767_en & bram_7_T_767_mask) begin
      bram_7[bram_7_T_767_addr] <= bram_7_T_767_data;
    end
    if(reset) begin
      state <= 2'h0;
    end else begin
      if(T_511) begin
        state <= 2'h0;
      end else begin
        if(T_504) begin
          if(T_502) begin
            state <= 2'h3;
          end else begin
            if(T_494) begin
              if(T_502) begin
                state <= 2'h0;
              end else begin
                if(T_482) begin
                  if(is_putblk) begin
                    state <= 2'h2;
                  end else begin
                    if(is_getblk) begin
                      state <= 2'h1;
                    end else begin
                      if(T_490) begin
                        state <= 2'h3;
                      end
                    end
                  end
                end
              end
            end else begin
              if(T_482) begin
                if(is_putblk) begin
                  state <= 2'h2;
                end else begin
                  if(is_getblk) begin
                    state <= 2'h1;
                  end else begin
                    if(T_490) begin
                      state <= 2'h3;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if(T_494) begin
            if(T_502) begin
              state <= 2'h0;
            end else begin
              if(T_482) begin
                if(is_putblk) begin
                  state <= 2'h2;
                end else begin
                  if(is_getblk) begin
                    state <= 2'h1;
                  end else begin
                    if(T_490) begin
                      state <= 2'h3;
                    end
                  end
                end
              end
            end
          end else begin
            if(T_482) begin
              if(is_putblk) begin
                state <= 2'h2;
              end else begin
                if(is_getblk) begin
                  state <= 2'h1;
                end else begin
                  if(T_490) begin
                    state <= 2'h3;
                  end
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_482) begin
        r_acq_addr_block <= io_acquire_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_482) begin
        r_acq_client_xact_id <= io_acquire_bits_client_xact_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_494) begin
        r_acq_addr_beat <= T_497;
      end else begin
        if(T_482) begin
          r_acq_addr_beat <= io_acquire_bits_addr_beat;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_482) begin
        r_acq_is_builtin_type <= io_acquire_bits_is_builtin_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_482) begin
        r_acq_a_type <= io_acquire_bits_a_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_482) begin
        r_acq_union <= io_acquire_bits_union;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_504) begin
        beats <= T_500;
      end else begin
        if(T_494) begin
          beats <= T_500;
        end else begin
          if(T_482) begin
            if(is_putblk) begin
              beats <= 3'h6;
            end else begin
              if(is_getblk) begin
                beats <= 3'h7;
              end
            end
          end
        end
      end
    end
  end
endmodule
module ReorderQueue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_data_addr_beat,
  input   io_enq_bits_data_subblock,
  input  [4:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [4:0] io_deq_tag,
  output [2:0] io_deq_data_addr_beat,
  output  io_deq_data_subblock,
  output  io_deq_matches
);
  reg [2:0] roq_data_addr_beat [0:3];
  reg [31:0] GEN_11;
  wire [2:0] roq_data_addr_beat_T_254_data;
  wire [1:0] roq_data_addr_beat_T_254_addr;
  wire  roq_data_addr_beat_T_254_en;
  wire [2:0] roq_data_addr_beat_T_276_data;
  wire [1:0] roq_data_addr_beat_T_276_addr;
  wire  roq_data_addr_beat_T_276_mask;
  wire  roq_data_addr_beat_T_276_en;
  reg  roq_data_subblock [0:3];
  reg [31:0] GEN_12;
  wire  roq_data_subblock_T_254_data;
  wire [1:0] roq_data_subblock_T_254_addr;
  wire  roq_data_subblock_T_254_en;
  wire  roq_data_subblock_T_276_data;
  wire [1:0] roq_data_subblock_T_276_addr;
  wire  roq_data_subblock_T_276_mask;
  wire  roq_data_subblock_T_276_en;
  reg [4:0] roq_tags_0;
  reg [31:0] GEN_13;
  reg [4:0] roq_tags_1;
  reg [31:0] GEN_14;
  reg [4:0] roq_tags_2;
  reg [31:0] GEN_15;
  reg [4:0] roq_tags_3;
  reg [31:0] GEN_16;
  wire  T_218_0;
  wire  T_218_1;
  wire  T_218_2;
  wire  T_218_3;
  reg  roq_free_0;
  reg [31:0] GEN_17;
  reg  roq_free_1;
  reg [31:0] GEN_18;
  reg  roq_free_2;
  reg [31:0] GEN_23;
  reg  roq_free_3;
  reg [31:0] GEN_32;
  wire [1:0] T_227;
  wire [1:0] T_228;
  wire [1:0] roq_enq_addr;
  wire  T_229;
  wire  T_231;
  wire  T_232;
  wire  T_233;
  wire  T_235;
  wire  T_236;
  wire  T_237;
  wire  T_239;
  wire  T_240;
  wire  T_241;
  wire  T_243;
  wire  T_244;
  wire [1:0] T_249;
  wire [1:0] T_250;
  wire [1:0] roq_deq_addr;
  wire  T_251;
  wire  T_252;
  wire  T_253;
  wire  T_272;
  wire  T_273;
  wire  T_274;
  wire  T_275;
  wire [4:0] GEN_0;
  wire [1:0] GEN_37;
  wire [4:0] GEN_3;
  wire [1:0] GEN_38;
  wire [4:0] GEN_4;
  wire [4:0] GEN_5;
  wire [4:0] GEN_6;
  wire  GEN_1;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [4:0] GEN_19;
  wire [4:0] GEN_20;
  wire [4:0] GEN_21;
  wire [4:0] GEN_22;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_2;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  assign io_enq_ready = T_253;
  assign io_deq_data_addr_beat = roq_data_addr_beat_T_254_data;
  assign io_deq_data_subblock = roq_data_subblock_T_254_data;
  assign io_deq_matches = T_274;
  assign roq_data_addr_beat_T_254_addr = roq_deq_addr;
  assign roq_data_addr_beat_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_addr_beat_T_254_data = roq_data_addr_beat[roq_data_addr_beat_T_254_addr];
  `else
  assign roq_data_addr_beat_T_254_data = roq_data_addr_beat_T_254_addr >= 3'h4 ? $random : roq_data_addr_beat[roq_data_addr_beat_T_254_addr];
  `endif
  assign roq_data_addr_beat_T_276_data = io_enq_bits_data_addr_beat;
  assign roq_data_addr_beat_T_276_addr = roq_enq_addr;
  assign roq_data_addr_beat_T_276_mask = T_275;
  assign roq_data_addr_beat_T_276_en = T_275;
  assign roq_data_subblock_T_254_addr = roq_deq_addr;
  assign roq_data_subblock_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_subblock_T_254_data = roq_data_subblock[roq_data_subblock_T_254_addr];
  `else
  assign roq_data_subblock_T_254_data = roq_data_subblock_T_254_addr >= 3'h4 ? $random : roq_data_subblock[roq_data_subblock_T_254_addr];
  `endif
  assign roq_data_subblock_T_276_data = io_enq_bits_data_subblock;
  assign roq_data_subblock_T_276_addr = roq_enq_addr;
  assign roq_data_subblock_T_276_mask = T_275;
  assign roq_data_subblock_T_276_en = T_275;
  assign T_218_0 = 1'h1;
  assign T_218_1 = 1'h1;
  assign T_218_2 = 1'h1;
  assign T_218_3 = 1'h1;
  assign T_227 = roq_free_2 ? 2'h2 : 2'h3;
  assign T_228 = roq_free_1 ? {{1'd0}, 1'h1} : T_227;
  assign roq_enq_addr = roq_free_0 ? {{1'd0}, 1'h0} : T_228;
  assign T_229 = roq_tags_0 == io_deq_tag;
  assign T_231 = roq_free_0 == 1'h0;
  assign T_232 = T_229 & T_231;
  assign T_233 = roq_tags_1 == io_deq_tag;
  assign T_235 = roq_free_1 == 1'h0;
  assign T_236 = T_233 & T_235;
  assign T_237 = roq_tags_2 == io_deq_tag;
  assign T_239 = roq_free_2 == 1'h0;
  assign T_240 = T_237 & T_239;
  assign T_241 = roq_tags_3 == io_deq_tag;
  assign T_243 = roq_free_3 == 1'h0;
  assign T_244 = T_241 & T_243;
  assign T_249 = T_240 ? 2'h2 : 2'h3;
  assign T_250 = T_236 ? {{1'd0}, 1'h1} : T_249;
  assign roq_deq_addr = T_232 ? {{1'd0}, 1'h0} : T_250;
  assign T_251 = roq_free_0 | roq_free_1;
  assign T_252 = T_251 | roq_free_2;
  assign T_253 = T_252 | roq_free_3;
  assign T_272 = T_232 | T_236;
  assign T_273 = T_272 | T_240;
  assign T_274 = T_273 | T_244;
  assign T_275 = io_enq_valid & io_enq_ready;
  assign GEN_0 = io_enq_bits_tag;
  assign GEN_37 = {{1'd0}, 1'h0};
  assign GEN_3 = GEN_37 == roq_enq_addr ? GEN_0 : roq_tags_0;
  assign GEN_38 = {{1'd0}, 1'h1};
  assign GEN_4 = GEN_38 == roq_enq_addr ? GEN_0 : roq_tags_1;
  assign GEN_5 = 2'h2 == roq_enq_addr ? GEN_0 : roq_tags_2;
  assign GEN_6 = 2'h3 == roq_enq_addr ? GEN_0 : roq_tags_3;
  assign GEN_1 = 1'h0;
  assign GEN_7 = GEN_37 == roq_enq_addr ? GEN_1 : roq_free_0;
  assign GEN_8 = GEN_38 == roq_enq_addr ? GEN_1 : roq_free_1;
  assign GEN_9 = 2'h2 == roq_enq_addr ? GEN_1 : roq_free_2;
  assign GEN_10 = 2'h3 == roq_enq_addr ? GEN_1 : roq_free_3;
  assign GEN_19 = T_275 ? GEN_3 : roq_tags_0;
  assign GEN_20 = T_275 ? GEN_4 : roq_tags_1;
  assign GEN_21 = T_275 ? GEN_5 : roq_tags_2;
  assign GEN_22 = T_275 ? GEN_6 : roq_tags_3;
  assign GEN_24 = T_275 ? GEN_7 : roq_free_0;
  assign GEN_25 = T_275 ? GEN_8 : roq_free_1;
  assign GEN_26 = T_275 ? GEN_9 : roq_free_2;
  assign GEN_27 = T_275 ? GEN_10 : roq_free_3;
  assign GEN_2 = 1'h1;
  assign GEN_28 = GEN_37 == roq_deq_addr ? GEN_2 : GEN_24;
  assign GEN_29 = GEN_38 == roq_deq_addr ? GEN_2 : GEN_25;
  assign GEN_30 = 2'h2 == roq_deq_addr ? GEN_2 : GEN_26;
  assign GEN_31 = 2'h3 == roq_deq_addr ? GEN_2 : GEN_27;
  assign GEN_33 = io_deq_valid ? GEN_28 : GEN_24;
  assign GEN_34 = io_deq_valid ? GEN_29 : GEN_25;
  assign GEN_35 = io_deq_valid ? GEN_30 : GEN_26;
  assign GEN_36 = io_deq_valid ? GEN_31 : GEN_27;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_11 = {1{$random}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    roq_data_addr_beat[initvar] = GEN_11[2:0];
  GEN_12 = {1{$random}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    roq_data_subblock[initvar] = GEN_12[0:0];
  GEN_13 = {1{$random}};
  roq_tags_0 = GEN_13[4:0];
  GEN_14 = {1{$random}};
  roq_tags_1 = GEN_14[4:0];
  GEN_15 = {1{$random}};
  roq_tags_2 = GEN_15[4:0];
  GEN_16 = {1{$random}};
  roq_tags_3 = GEN_16[4:0];
  GEN_17 = {1{$random}};
  roq_free_0 = GEN_17[0:0];
  GEN_18 = {1{$random}};
  roq_free_1 = GEN_18[0:0];
  GEN_23 = {1{$random}};
  roq_free_2 = GEN_23[0:0];
  GEN_32 = {1{$random}};
  roq_free_3 = GEN_32[0:0];
  end
`endif
  always @(posedge clk) begin
    if(roq_data_addr_beat_T_276_en & roq_data_addr_beat_T_276_mask) begin
      roq_data_addr_beat[roq_data_addr_beat_T_276_addr] <= roq_data_addr_beat_T_276_data;
    end
    if(roq_data_subblock_T_276_en & roq_data_subblock_T_276_mask) begin
      roq_data_subblock[roq_data_subblock_T_276_addr] <= roq_data_subblock_T_276_data;
    end
    if(1'h0) begin
    end else begin
      if(T_275) begin
        if(GEN_37 == roq_enq_addr) begin
          roq_tags_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_275) begin
        if(GEN_38 == roq_enq_addr) begin
          roq_tags_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_275) begin
        if(2'h2 == roq_enq_addr) begin
          roq_tags_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_275) begin
        if(2'h3 == roq_enq_addr) begin
          roq_tags_3 <= GEN_0;
        end
      end
    end
    if(reset) begin
      roq_free_0 <= T_218_0;
    end else begin
      if(io_deq_valid) begin
        if(GEN_37 == roq_deq_addr) begin
          roq_free_0 <= GEN_2;
        end else begin
          if(T_275) begin
            if(GEN_37 == roq_enq_addr) begin
              roq_free_0 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_275) begin
          if(GEN_37 == roq_enq_addr) begin
            roq_free_0 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_1 <= T_218_1;
    end else begin
      if(io_deq_valid) begin
        if(GEN_38 == roq_deq_addr) begin
          roq_free_1 <= GEN_2;
        end else begin
          if(T_275) begin
            if(GEN_38 == roq_enq_addr) begin
              roq_free_1 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_275) begin
          if(GEN_38 == roq_enq_addr) begin
            roq_free_1 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_2 <= T_218_2;
    end else begin
      if(io_deq_valid) begin
        if(2'h2 == roq_deq_addr) begin
          roq_free_2 <= GEN_2;
        end else begin
          if(T_275) begin
            if(2'h2 == roq_enq_addr) begin
              roq_free_2 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_275) begin
          if(2'h2 == roq_enq_addr) begin
            roq_free_2 <= GEN_1;
          end
        end
      end
    end
    if(reset) begin
      roq_free_3 <= T_218_3;
    end else begin
      if(io_deq_valid) begin
        if(2'h3 == roq_deq_addr) begin
          roq_free_3 <= GEN_2;
        end else begin
          if(T_275) begin
            if(2'h3 == roq_enq_addr) begin
              roq_free_3 <= GEN_1;
            end
          end
        end
      end else begin
        if(T_275) begin
          if(2'h3 == roq_enq_addr) begin
            roq_free_3 <= GEN_1;
          end
        end
      end
    end
  end
endmodule
module NastiIOTileLinkIOIdMapper_2(
  input   clk,
  input   reset,
  input   io_req_valid,
  output  io_req_ready,
  input  [1:0] io_req_tl_id,
  output [4:0] io_req_nasti_id,
  input   io_resp_valid,
  output  io_resp_matches,
  input  [4:0] io_resp_nasti_id,
  output [1:0] io_resp_tl_id
);
  assign io_req_ready = 1'h1;
  assign io_req_nasti_id = {{3'd0}, io_req_tl_id};
  assign io_resp_matches = 1'h1;
  assign io_resp_tl_id = io_resp_nasti_id[1:0];
endmodule
module Arbiter_14(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output  io_chosen
);
  wire  GEN_0;
  wire [2:0] GEN_1;
  wire [1:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire [3:0] GEN_5;
  wire [63:0] GEN_6;
  wire  GEN_7;
  wire  T_542;
  wire  T_544;
  wire  T_546;
  wire  T_547;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_544;
  assign io_out_valid = T_547;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_client_id = GEN_7;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr_beat : io_in_1_bits_addr_beat;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_client_xact_id : io_in_1_bits_client_xact_id;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_manager_xact_id : io_in_1_bits_manager_xact_id;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_is_builtin_type : io_in_1_bits_is_builtin_type;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_g_type : io_in_1_bits_g_type;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_client_id : io_in_1_bits_client_id;
  assign T_542 = io_in_0_valid == 1'h0;
  assign T_544 = T_542 & io_out_ready;
  assign T_546 = T_542 == 1'h0;
  assign T_547 = T_546 | io_in_1_valid;
endmodule
module NastiIOTileLinkIOConverter_1(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  input   io_nasti_aw_ready,
  output  io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  output [7:0] io_nasti_aw_bits_len,
  output [2:0] io_nasti_aw_bits_size,
  output [1:0] io_nasti_aw_bits_burst,
  output  io_nasti_aw_bits_lock,
  output [3:0] io_nasti_aw_bits_cache,
  output [2:0] io_nasti_aw_bits_prot,
  output [3:0] io_nasti_aw_bits_qos,
  output [3:0] io_nasti_aw_bits_region,
  output [4:0] io_nasti_aw_bits_id,
  output  io_nasti_aw_bits_user,
  input   io_nasti_w_ready,
  output  io_nasti_w_valid,
  output [63:0] io_nasti_w_bits_data,
  output  io_nasti_w_bits_last,
  output [4:0] io_nasti_w_bits_id,
  output [7:0] io_nasti_w_bits_strb,
  output  io_nasti_w_bits_user,
  output  io_nasti_b_ready,
  input   io_nasti_b_valid,
  input  [1:0] io_nasti_b_bits_resp,
  input  [4:0] io_nasti_b_bits_id,
  input   io_nasti_b_bits_user,
  input   io_nasti_ar_ready,
  output  io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output [7:0] io_nasti_ar_bits_len,
  output [2:0] io_nasti_ar_bits_size,
  output [1:0] io_nasti_ar_bits_burst,
  output  io_nasti_ar_bits_lock,
  output [3:0] io_nasti_ar_bits_cache,
  output [2:0] io_nasti_ar_bits_prot,
  output [3:0] io_nasti_ar_bits_qos,
  output [3:0] io_nasti_ar_bits_region,
  output [4:0] io_nasti_ar_bits_id,
  output  io_nasti_ar_bits_user,
  output  io_nasti_r_ready,
  input   io_nasti_r_valid,
  input  [1:0] io_nasti_r_bits_resp,
  input  [63:0] io_nasti_r_bits_data,
  input   io_nasti_r_bits_last,
  input  [4:0] io_nasti_r_bits_id,
  input   io_nasti_r_bits_user
);
  wire [2:0] T_593_0;
  wire [2:0] T_593_1;
  wire [2:0] T_593_2;
  wire  T_595;
  wire  T_596;
  wire  T_597;
  wire  T_600;
  wire  T_601;
  wire  has_data;
  wire [2:0] T_610_0;
  wire [2:0] T_610_1;
  wire [2:0] T_610_2;
  wire  T_612;
  wire  T_613;
  wire  T_614;
  wire  T_617;
  wire  T_618;
  wire  is_subblock;
  wire [2:0] T_627_0;
  wire  T_629;
  wire  is_multibeat;
  wire  T_632;
  wire  T_633;
  reg [2:0] tl_cnt_out;
  reg [31:0] GEN_15;
  wire  T_636;
  wire [2:0] GEN_6;
  wire [3:0] T_638;
  wire [2:0] T_639;
  wire [2:0] GEN_0;
  wire  tl_wrap_out;
  wire  T_641;
  wire  get_valid;
  wire  put_valid;
  wire  roq_clk;
  wire  roq_reset;
  wire  roq_io_enq_ready;
  wire  roq_io_enq_valid;
  wire [2:0] roq_io_enq_bits_data_addr_beat;
  wire  roq_io_enq_bits_data_subblock;
  wire [4:0] roq_io_enq_bits_tag;
  wire  roq_io_deq_valid;
  wire [4:0] roq_io_deq_tag;
  wire [2:0] roq_io_deq_data_addr_beat;
  wire  roq_io_deq_data_subblock;
  wire  roq_io_deq_matches;
  wire  get_id_mapper_clk;
  wire  get_id_mapper_reset;
  wire  get_id_mapper_io_req_valid;
  wire  get_id_mapper_io_req_ready;
  wire [1:0] get_id_mapper_io_req_tl_id;
  wire [4:0] get_id_mapper_io_req_nasti_id;
  wire  get_id_mapper_io_resp_valid;
  wire  get_id_mapper_io_resp_matches;
  wire [4:0] get_id_mapper_io_resp_nasti_id;
  wire [1:0] get_id_mapper_io_resp_tl_id;
  wire  put_id_mapper_clk;
  wire  put_id_mapper_reset;
  wire  put_id_mapper_io_req_valid;
  wire  put_id_mapper_io_req_ready;
  wire [1:0] put_id_mapper_io_req_tl_id;
  wire [4:0] put_id_mapper_io_req_nasti_id;
  wire  put_id_mapper_io_resp_valid;
  wire  put_id_mapper_io_resp_matches;
  wire [4:0] put_id_mapper_io_resp_nasti_id;
  wire [1:0] put_id_mapper_io_resp_tl_id;
  wire [2:0] GEN_7;
  wire  T_661;
  wire  put_id_mask;
  wire  T_663;
  wire  put_id_ready;
  reg  w_inflight;
  reg [31:0] GEN_16;
  wire  aw_ready;
  wire  T_665;
  wire  T_667;
  wire  T_668;
  reg [2:0] nasti_cnt_out;
  reg [31:0] GEN_17;
  wire  T_671;
  wire [3:0] T_673;
  wire [2:0] T_674;
  wire [2:0] GEN_1;
  wire  nasti_wrap_out;
  wire  T_675;
  wire  T_676;
  wire  T_678;
  wire  T_679;
  wire  T_680;
  wire  T_681;
  wire  T_683;
  wire  T_684;
  wire  T_685;
  wire  T_686;
  wire  T_687;
  wire  T_689;
  wire [2:0] T_690;
  wire [28:0] T_691;
  wire [31:0] T_692;
  wire [2:0] T_693;
  wire  T_703;
  wire [2:0] T_704;
  wire  T_705;
  wire [2:0] T_706;
  wire  T_707;
  wire [2:0] T_708;
  wire  T_709;
  wire [2:0] T_710;
  wire  T_711;
  wire [2:0] T_712;
  wire  T_713;
  wire [2:0] T_714;
  wire  T_715;
  wire [2:0] T_716;
  wire  T_717;
  wire [2:0] T_718;
  wire [2:0] T_720;
  wire [2:0] T_723;
  wire [31:0] T_736_addr;
  wire [7:0] T_736_len;
  wire [2:0] T_736_size;
  wire [1:0] T_736_burst;
  wire  T_736_lock;
  wire [3:0] T_736_cache;
  wire [2:0] T_736_prot;
  wire [3:0] T_736_qos;
  wire [3:0] T_736_region;
  wire [4:0] T_736_id;
  wire  T_736_user;
  wire  T_755;
  wire  T_756;
  wire  T_757;
  wire  T_758;
  wire [2:0] T_765;
  wire [31:0] T_778_addr;
  wire [7:0] T_778_len;
  wire [2:0] T_778_size;
  wire [1:0] T_778_burst;
  wire  T_778_lock;
  wire [3:0] T_778_cache;
  wire [2:0] T_778_prot;
  wire [3:0] T_778_qos;
  wire [3:0] T_778_region;
  wire [4:0] T_778_id;
  wire  T_778_user;
  wire  T_797;
  wire  T_799;
  wire  T_800;
  wire [7:0] GEN_9;
  wire [8:0] T_804;
  wire [7:0] T_805;
  wire [7:0] T_811_0;
  wire  T_814;
  wire  T_815;
  wire  T_817;
  wire  T_818;
  wire  T_819;
  wire [7:0] T_820;
  wire [7:0] T_822;
  wire [7:0] T_823;
  wire  T_825;
  wire  T_826;
  wire [63:0] T_833_data;
  wire  T_833_last;
  wire [4:0] T_833_id;
  wire [7:0] T_833_strb;
  wire  T_833_user;
  wire  T_844;
  wire  T_845;
  wire  T_846;
  wire  T_847;
  wire  T_848;
  wire  T_852;
  wire  T_853;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  T_856;
  wire [2:0] T_864_0;
  wire [3:0] GEN_10;
  wire  T_866;
  wire  T_874_0;
  wire [3:0] GEN_11;
  wire  T_876;
  wire  T_879;
  wire  T_881;
  reg [2:0] tl_cnt_in;
  reg [31:0] GEN_18;
  wire [3:0] T_886;
  wire [2:0] T_887;
  wire [2:0] GEN_5;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_0_bits_client_id;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_1_bits_client_id;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_out_bits_client_id;
  wire  gnt_arb_io_chosen;
  wire [2:0] T_914;
  wire [2:0] T_916;
  wire [2:0] T_939_addr_beat;
  wire [1:0] T_939_client_xact_id;
  wire  T_939_manager_xact_id;
  wire  T_939_is_builtin_type;
  wire [3:0] T_939_g_type;
  wire [63:0] T_939_data;
  wire  T_962;
  wire  T_963;
  wire  T_964;
  wire  T_966;
  wire  T_968;
  wire  T_969;
  wire  T_970;
  wire  T_972;
  wire [2:0] T_1000_addr_beat;
  wire [1:0] T_1000_client_xact_id;
  wire  T_1000_manager_xact_id;
  wire  T_1000_is_builtin_type;
  wire [3:0] T_1000_g_type;
  wire [63:0] T_1000_data;
  wire  T_1023;
  wire  T_1024;
  wire  T_1025;
  wire  T_1027;
  wire  T_1029;
  wire [1:0] GEN_13;
  wire  T_1031;
  wire  T_1032;
  wire  T_1033;
  wire  T_1035;
  wire  T_1037;
  wire  T_1039;
  wire  T_1040;
  wire  T_1041;
  wire  T_1043;
  reg [4:0] GEN_8;
  reg [31:0] GEN_19;
  reg  GEN_12;
  reg [31:0] GEN_20;
  reg  GEN_14;
  reg [31:0] GEN_21;
  ReorderQueue_3 roq (
    .clk(roq_clk),
    .reset(roq_reset),
    .io_enq_ready(roq_io_enq_ready),
    .io_enq_valid(roq_io_enq_valid),
    .io_enq_bits_data_addr_beat(roq_io_enq_bits_data_addr_beat),
    .io_enq_bits_data_subblock(roq_io_enq_bits_data_subblock),
    .io_enq_bits_tag(roq_io_enq_bits_tag),
    .io_deq_valid(roq_io_deq_valid),
    .io_deq_tag(roq_io_deq_tag),
    .io_deq_data_addr_beat(roq_io_deq_data_addr_beat),
    .io_deq_data_subblock(roq_io_deq_data_subblock),
    .io_deq_matches(roq_io_deq_matches)
  );
  NastiIOTileLinkIOIdMapper_2 get_id_mapper (
    .clk(get_id_mapper_clk),
    .reset(get_id_mapper_reset),
    .io_req_valid(get_id_mapper_io_req_valid),
    .io_req_ready(get_id_mapper_io_req_ready),
    .io_req_tl_id(get_id_mapper_io_req_tl_id),
    .io_req_nasti_id(get_id_mapper_io_req_nasti_id),
    .io_resp_valid(get_id_mapper_io_resp_valid),
    .io_resp_matches(get_id_mapper_io_resp_matches),
    .io_resp_nasti_id(get_id_mapper_io_resp_nasti_id),
    .io_resp_tl_id(get_id_mapper_io_resp_tl_id)
  );
  NastiIOTileLinkIOIdMapper_2 put_id_mapper (
    .clk(put_id_mapper_clk),
    .reset(put_id_mapper_reset),
    .io_req_valid(put_id_mapper_io_req_valid),
    .io_req_ready(put_id_mapper_io_req_ready),
    .io_req_tl_id(put_id_mapper_io_req_tl_id),
    .io_req_nasti_id(put_id_mapper_io_req_nasti_id),
    .io_resp_valid(put_id_mapper_io_resp_valid),
    .io_resp_matches(put_id_mapper_io_resp_matches),
    .io_resp_nasti_id(put_id_mapper_io_resp_nasti_id),
    .io_resp_tl_id(put_id_mapper_io_resp_tl_id)
  );
  Arbiter_14 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_0_bits_client_id(gnt_arb_io_in_0_bits_client_id),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_1_bits_client_id(gnt_arb_io_in_1_bits_client_id),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_out_bits_client_id(gnt_arb_io_out_bits_client_id),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_tl_acquire_ready = T_848;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_nasti_aw_valid = T_758;
  assign io_nasti_aw_bits_addr = T_778_addr;
  assign io_nasti_aw_bits_len = T_778_len;
  assign io_nasti_aw_bits_size = T_778_size;
  assign io_nasti_aw_bits_burst = T_778_burst;
  assign io_nasti_aw_bits_lock = T_778_lock;
  assign io_nasti_aw_bits_cache = T_778_cache;
  assign io_nasti_aw_bits_prot = T_778_prot;
  assign io_nasti_aw_bits_qos = T_778_qos;
  assign io_nasti_aw_bits_region = T_778_region;
  assign io_nasti_aw_bits_id = T_778_id;
  assign io_nasti_aw_bits_user = T_778_user;
  assign io_nasti_w_valid = T_797;
  assign io_nasti_w_bits_data = T_833_data;
  assign io_nasti_w_bits_last = T_833_last;
  assign io_nasti_w_bits_id = T_833_id;
  assign io_nasti_w_bits_strb = T_833_strb;
  assign io_nasti_w_bits_user = T_833_user;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_ar_valid = T_689;
  assign io_nasti_ar_bits_addr = T_736_addr;
  assign io_nasti_ar_bits_len = T_736_len;
  assign io_nasti_ar_bits_size = T_736_size;
  assign io_nasti_ar_bits_burst = T_736_burst;
  assign io_nasti_ar_bits_lock = T_736_lock;
  assign io_nasti_ar_bits_cache = T_736_cache;
  assign io_nasti_ar_bits_prot = T_736_prot;
  assign io_nasti_ar_bits_qos = T_736_qos;
  assign io_nasti_ar_bits_region = T_736_region;
  assign io_nasti_ar_bits_id = T_736_id;
  assign io_nasti_ar_bits_user = T_736_user;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign T_593_0 = 3'h2;
  assign T_593_1 = 3'h3;
  assign T_593_2 = 3'h4;
  assign T_595 = T_593_0 == io_tl_acquire_bits_a_type;
  assign T_596 = T_593_1 == io_tl_acquire_bits_a_type;
  assign T_597 = T_593_2 == io_tl_acquire_bits_a_type;
  assign T_600 = T_595 | T_596;
  assign T_601 = T_600 | T_597;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T_601;
  assign T_610_0 = 3'h2;
  assign T_610_1 = 3'h0;
  assign T_610_2 = 3'h4;
  assign T_612 = T_610_0 == io_tl_acquire_bits_a_type;
  assign T_613 = T_610_1 == io_tl_acquire_bits_a_type;
  assign T_614 = T_610_2 == io_tl_acquire_bits_a_type;
  assign T_617 = T_612 | T_613;
  assign T_618 = T_617 | T_614;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T_618;
  assign T_627_0 = 3'h3;
  assign T_629 = T_627_0 == io_tl_acquire_bits_a_type;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T_629;
  assign T_632 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T_633 = T_632 & is_multibeat;
  assign T_636 = tl_cnt_out == 3'h7;
  assign GEN_6 = {{2'd0}, 1'h1};
  assign T_638 = tl_cnt_out + GEN_6;
  assign T_639 = T_638[2:0];
  assign GEN_0 = T_633 ? T_639 : tl_cnt_out;
  assign tl_wrap_out = T_633 & T_636;
  assign T_641 = has_data == 1'h0;
  assign get_valid = io_tl_acquire_valid & T_641;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign roq_clk = clk;
  assign roq_reset = reset;
  assign roq_io_enq_valid = T_676;
  assign roq_io_enq_bits_data_addr_beat = io_tl_acquire_bits_addr_beat;
  assign roq_io_enq_bits_data_subblock = is_subblock;
  assign roq_io_enq_bits_tag = io_nasti_ar_bits_id;
  assign roq_io_deq_valid = T_679;
  assign roq_io_deq_tag = io_nasti_r_bits_id;
  assign get_id_mapper_clk = clk;
  assign get_id_mapper_reset = reset;
  assign get_id_mapper_io_req_valid = T_681;
  assign get_id_mapper_io_req_tl_id = io_tl_acquire_bits_client_xact_id;
  assign get_id_mapper_io_resp_valid = T_683;
  assign get_id_mapper_io_resp_nasti_id = io_nasti_r_bits_id;
  assign put_id_mapper_clk = clk;
  assign put_id_mapper_reset = reset;
  assign put_id_mapper_io_req_valid = T_686;
  assign put_id_mapper_io_req_tl_id = io_tl_acquire_bits_client_xact_id;
  assign put_id_mapper_io_resp_valid = T_687;
  assign put_id_mapper_io_resp_nasti_id = io_nasti_b_bits_id;
  assign GEN_7 = {{2'd0}, 1'h0};
  assign T_661 = io_tl_acquire_bits_addr_beat == GEN_7;
  assign put_id_mask = is_subblock | T_661;
  assign T_663 = put_id_mask == 1'h0;
  assign put_id_ready = put_id_mapper_io_req_ready | T_663;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T_665 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_667 = roq_io_deq_data_subblock == 1'h0;
  assign T_668 = T_665 & T_667;
  assign T_671 = nasti_cnt_out == 3'h7;
  assign T_673 = nasti_cnt_out + GEN_6;
  assign T_674 = T_673[2:0];
  assign GEN_1 = T_668 ? T_674 : nasti_cnt_out;
  assign nasti_wrap_out = T_668 & T_671;
  assign T_675 = get_valid & io_nasti_ar_ready;
  assign T_676 = T_675 & get_id_mapper_io_req_ready;
  assign T_678 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign T_679 = T_665 & T_678;
  assign T_680 = get_valid & roq_io_enq_ready;
  assign T_681 = T_680 & io_nasti_ar_ready;
  assign T_683 = T_665 & io_nasti_r_bits_last;
  assign T_684 = put_valid & aw_ready;
  assign T_685 = T_684 & io_nasti_w_ready;
  assign T_686 = T_685 & put_id_mask;
  assign T_687 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_689 = T_680 & get_id_mapper_io_req_ready;
  assign T_690 = io_tl_acquire_bits_union[11:9];
  assign T_691 = {io_tl_acquire_bits_addr_block,io_tl_acquire_bits_addr_beat};
  assign T_692 = {T_691,T_690};
  assign T_693 = io_tl_acquire_bits_union[8:6];
  assign T_703 = 3'h7 == T_693;
  assign T_704 = T_703 ? {{1'd0}, 2'h3} : 3'h7;
  assign T_705 = 3'h3 == T_693;
  assign T_706 = T_705 ? {{1'd0}, 2'h3} : T_704;
  assign T_707 = 3'h6 == T_693;
  assign T_708 = T_707 ? {{1'd0}, 2'h2} : T_706;
  assign T_709 = 3'h2 == T_693;
  assign T_710 = T_709 ? {{1'd0}, 2'h2} : T_708;
  assign T_711 = 3'h5 == T_693;
  assign T_712 = T_711 ? {{2'd0}, 1'h1} : T_710;
  assign T_713 = 3'h1 == T_693;
  assign T_714 = T_713 ? {{2'd0}, 1'h1} : T_712;
  assign T_715 = 3'h4 == T_693;
  assign T_716 = T_715 ? {{2'd0}, 1'h0} : T_714;
  assign T_717 = 3'h0 == T_693;
  assign T_718 = T_717 ? {{2'd0}, 1'h0} : T_716;
  assign T_720 = is_subblock ? T_718 : {{1'd0}, 2'h3};
  assign T_723 = is_subblock ? {{2'd0}, 1'h0} : 3'h7;
  assign T_736_addr = T_692;
  assign T_736_len = {{5'd0}, T_723};
  assign T_736_size = T_720;
  assign T_736_burst = 2'h1;
  assign T_736_lock = 1'h0;
  assign T_736_cache = {{3'd0}, 1'h0};
  assign T_736_prot = {{2'd0}, 1'h0};
  assign T_736_qos = {{3'd0}, 1'h0};
  assign T_736_region = {{3'd0}, 1'h0};
  assign T_736_id = get_id_mapper_io_req_nasti_id;
  assign T_736_user = 1'h0;
  assign T_755 = w_inflight == 1'h0;
  assign T_756 = put_valid & io_nasti_w_ready;
  assign T_757 = T_756 & put_id_ready;
  assign T_758 = T_757 & T_755;
  assign T_765 = is_multibeat ? 3'h7 : {{2'd0}, 1'h0};
  assign T_778_addr = T_692;
  assign T_778_len = {{5'd0}, T_765};
  assign T_778_size = {{1'd0}, 2'h3};
  assign T_778_burst = 2'h1;
  assign T_778_lock = 1'h0;
  assign T_778_cache = 4'h0;
  assign T_778_prot = 3'h0;
  assign T_778_qos = 4'h0;
  assign T_778_region = 4'h0;
  assign T_778_id = put_id_mapper_io_req_nasti_id;
  assign T_778_user = 1'h0;
  assign T_797 = T_684 & put_id_ready;
  assign T_799 = io_tl_acquire_bits_a_type == 3'h4;
  assign T_800 = io_tl_acquire_bits_is_builtin_type & T_799;
  assign GEN_9 = {{7'd0}, 1'h1};
  assign T_804 = 8'h0 - GEN_9;
  assign T_805 = T_804[7:0];
  assign T_811_0 = T_805;
  assign T_814 = io_tl_acquire_bits_a_type == 3'h3;
  assign T_815 = io_tl_acquire_bits_is_builtin_type & T_814;
  assign T_817 = io_tl_acquire_bits_a_type == 3'h2;
  assign T_818 = io_tl_acquire_bits_is_builtin_type & T_817;
  assign T_819 = T_815 | T_818;
  assign T_820 = io_tl_acquire_bits_union[8:1];
  assign T_822 = T_819 ? T_820 : {{7'd0}, 1'h0};
  assign T_823 = T_800 ? T_811_0 : T_822;
  assign T_825 = T_632 & is_subblock;
  assign T_826 = tl_wrap_out | T_825;
  assign T_833_data = io_tl_acquire_bits_data;
  assign T_833_last = T_826;
  assign T_833_id = GEN_8;
  assign T_833_strb = T_823;
  assign T_833_user = 1'h0;
  assign T_844 = aw_ready & io_nasti_w_ready;
  assign T_845 = T_844 & put_id_ready;
  assign T_846 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T_847 = T_846 & get_id_mapper_io_req_ready;
  assign T_848 = has_data ? T_845 : T_847;
  assign T_852 = T_755 & T_632;
  assign T_853 = T_852 & is_multibeat;
  assign GEN_2 = T_853 ? 1'h1 : w_inflight;
  assign GEN_3 = tl_wrap_out ? 1'h0 : GEN_2;
  assign GEN_4 = w_inflight ? GEN_3 : GEN_2;
  assign T_856 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_864_0 = 3'h5;
  assign GEN_10 = {{1'd0}, T_864_0};
  assign T_866 = GEN_10 == io_tl_grant_bits_g_type;
  assign T_874_0 = 1'h0;
  assign GEN_11 = {{3'd0}, T_874_0};
  assign T_876 = GEN_11 == io_tl_grant_bits_g_type;
  assign T_879 = io_tl_grant_bits_is_builtin_type ? T_866 : T_876;
  assign T_881 = T_856 & T_879;
  assign T_886 = tl_cnt_in + GEN_6;
  assign T_887 = T_886[2:0];
  assign GEN_5 = T_881 ? T_887 : tl_cnt_in;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_nasti_r_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = T_939_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = T_939_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = T_939_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = T_939_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = T_939_g_type;
  assign gnt_arb_io_in_0_bits_data = T_939_data;
  assign gnt_arb_io_in_0_bits_client_id = GEN_12;
  assign gnt_arb_io_in_1_valid = io_nasti_b_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = T_1000_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = T_1000_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = T_1000_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = T_1000_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = T_1000_g_type;
  assign gnt_arb_io_in_1_bits_data = T_1000_data;
  assign gnt_arb_io_in_1_bits_client_id = GEN_14;
  assign gnt_arb_io_out_ready = io_tl_grant_ready;
  assign T_914 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T_916 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T_939_addr_beat = T_916;
  assign T_939_client_xact_id = get_id_mapper_io_resp_tl_id;
  assign T_939_manager_xact_id = 1'h0;
  assign T_939_is_builtin_type = 1'h1;
  assign T_939_g_type = {{1'd0}, T_914};
  assign T_939_data = io_nasti_r_bits_data;
  assign T_962 = roq_io_deq_valid == 1'h0;
  assign T_963 = T_962 | roq_io_deq_matches;
  assign T_964 = T_963 | reset;
  assign T_966 = T_964 == 1'h0;
  assign T_968 = gnt_arb_io_in_0_valid == 1'h0;
  assign T_969 = T_968 | get_id_mapper_io_resp_matches;
  assign T_970 = T_969 | reset;
  assign T_972 = T_970 == 1'h0;
  assign T_1000_addr_beat = {{2'd0}, 1'h0};
  assign T_1000_client_xact_id = put_id_mapper_io_resp_tl_id;
  assign T_1000_manager_xact_id = 1'h0;
  assign T_1000_is_builtin_type = 1'h1;
  assign T_1000_g_type = {{1'd0}, 3'h3};
  assign T_1000_data = {{63'd0}, 1'h0};
  assign T_1023 = gnt_arb_io_in_1_valid == 1'h0;
  assign T_1024 = T_1023 | put_id_mapper_io_resp_matches;
  assign T_1025 = T_1024 | reset;
  assign T_1027 = T_1025 == 1'h0;
  assign T_1029 = io_nasti_r_valid == 1'h0;
  assign GEN_13 = {{1'd0}, 1'h0};
  assign T_1031 = io_nasti_r_bits_resp == GEN_13;
  assign T_1032 = T_1029 | T_1031;
  assign T_1033 = T_1032 | reset;
  assign T_1035 = T_1033 == 1'h0;
  assign T_1037 = io_nasti_b_valid == 1'h0;
  assign T_1039 = io_nasti_b_bits_resp == GEN_13;
  assign T_1040 = T_1037 | T_1039;
  assign T_1041 = T_1040 | reset;
  assign T_1043 = T_1041 == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  tl_cnt_out = GEN_15[2:0];
  GEN_16 = {1{$random}};
  w_inflight = GEN_16[0:0];
  GEN_17 = {1{$random}};
  nasti_cnt_out = GEN_17[2:0];
  GEN_18 = {1{$random}};
  tl_cnt_in = GEN_18[2:0];
  GEN_19 = {1{$random}};
  GEN_8 = GEN_19[4:0];
  GEN_20 = {1{$random}};
  GEN_12 = GEN_20[0:0];
  GEN_21 = {1{$random}};
  GEN_14 = GEN_21[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else begin
      if(T_633) begin
        tl_cnt_out <= T_639;
      end
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else begin
      if(w_inflight) begin
        if(tl_wrap_out) begin
          w_inflight <= 1'h0;
        end else begin
          if(T_853) begin
            w_inflight <= 1'h1;
          end
        end
      end else begin
        if(T_853) begin
          w_inflight <= 1'h1;
        end
      end
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else begin
      if(T_668) begin
        nasti_cnt_out <= T_674;
      end
    end
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else begin
      if(T_881) begin
        tl_cnt_in <= T_887;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_966) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI converter ReorderQueue: NASTI tag error\n    at Nasti.scala:210 assert(!roq.io.deq.valid || roq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_966) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_966) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_972) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI ID Mapper: NASTI tag error\n    at Nasti.scala:212 assert(!gnt_arb.io.in(0).valid || get_id_mapper.io.resp.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_972) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_972) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1027) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at Nasti.scala:224 assert(!gnt_arb.io.in(1).valid || put_id_mapper.io.resp.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1027) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1027) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1035) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI read error\n    at Nasti.scala:226 assert(!io.nasti.r.valid || io.nasti.r.bits.resp === UInt(0), \"NASTI read error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1035) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1035) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1043) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI write error\n    at Nasti.scala:227 assert(!io.nasti.b.valid || io.nasti.b.bits.resp === UInt(0), \"NASTI write error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1043) begin
          $fwrite(32'h80000002,"1\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1043) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Uncore(
  input   clk,
  input   reset,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  output  io_tiles_cached_0_acquire_ready,
  input   io_tiles_cached_0_acquire_valid,
  input  [25:0] io_tiles_cached_0_acquire_bits_addr_block,
  input  [1:0] io_tiles_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_cached_0_acquire_bits_addr_beat,
  input   io_tiles_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_cached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_cached_0_acquire_bits_union,
  input  [63:0] io_tiles_cached_0_acquire_bits_data,
  input   io_tiles_cached_0_probe_ready,
  output  io_tiles_cached_0_probe_valid,
  output [25:0] io_tiles_cached_0_probe_bits_addr_block,
  output [1:0] io_tiles_cached_0_probe_bits_p_type,
  output  io_tiles_cached_0_release_ready,
  input   io_tiles_cached_0_release_valid,
  input  [2:0] io_tiles_cached_0_release_bits_addr_beat,
  input  [25:0] io_tiles_cached_0_release_bits_addr_block,
  input  [1:0] io_tiles_cached_0_release_bits_client_xact_id,
  input   io_tiles_cached_0_release_bits_voluntary,
  input  [2:0] io_tiles_cached_0_release_bits_r_type,
  input  [63:0] io_tiles_cached_0_release_bits_data,
  input   io_tiles_cached_0_grant_ready,
  output  io_tiles_cached_0_grant_valid,
  output [2:0] io_tiles_cached_0_grant_bits_addr_beat,
  output [1:0] io_tiles_cached_0_grant_bits_client_xact_id,
  output [2:0] io_tiles_cached_0_grant_bits_manager_xact_id,
  output  io_tiles_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_cached_0_grant_bits_g_type,
  output [63:0] io_tiles_cached_0_grant_bits_data,
  output  io_tiles_cached_0_grant_bits_manager_id,
  output  io_tiles_cached_0_finish_ready,
  input   io_tiles_cached_0_finish_valid,
  input  [2:0] io_tiles_cached_0_finish_bits_manager_xact_id,
  input   io_tiles_cached_0_finish_bits_manager_id,
  output  io_tiles_uncached_0_acquire_ready,
  input   io_tiles_uncached_0_acquire_valid,
  input  [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
  input  [1:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_uncached_0_acquire_bits_addr_beat,
  input   io_tiles_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_uncached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_uncached_0_acquire_bits_union,
  input  [63:0] io_tiles_uncached_0_acquire_bits_data,
  input   io_tiles_uncached_0_grant_ready,
  output  io_tiles_uncached_0_grant_valid,
  output [2:0] io_tiles_uncached_0_grant_bits_addr_beat,
  output [1:0] io_tiles_uncached_0_grant_bits_client_xact_id,
  output [2:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
  output  io_tiles_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_uncached_0_grant_bits_g_type,
  output [63:0] io_tiles_uncached_0_grant_bits_data,
  output  io_prci_0_reset,
  output  io_prci_0_id,
  output  io_prci_0_interrupts_meip,
  output  io_prci_0_interrupts_seip,
  output  io_prci_0_interrupts_debug,
  output  io_prci_0_interrupts_mtip,
  output  io_prci_0_interrupts_msip,
  input   io_mmio_axi_0_aw_ready,
  output  io_mmio_axi_0_aw_valid,
  output [31:0] io_mmio_axi_0_aw_bits_addr,
  output [7:0] io_mmio_axi_0_aw_bits_len,
  output [2:0] io_mmio_axi_0_aw_bits_size,
  output [1:0] io_mmio_axi_0_aw_bits_burst,
  output  io_mmio_axi_0_aw_bits_lock,
  output [3:0] io_mmio_axi_0_aw_bits_cache,
  output [2:0] io_mmio_axi_0_aw_bits_prot,
  output [3:0] io_mmio_axi_0_aw_bits_qos,
  output [3:0] io_mmio_axi_0_aw_bits_region,
  output [4:0] io_mmio_axi_0_aw_bits_id,
  output  io_mmio_axi_0_aw_bits_user,
  input   io_mmio_axi_0_w_ready,
  output  io_mmio_axi_0_w_valid,
  output [63:0] io_mmio_axi_0_w_bits_data,
  output  io_mmio_axi_0_w_bits_last,
  output [4:0] io_mmio_axi_0_w_bits_id,
  output [7:0] io_mmio_axi_0_w_bits_strb,
  output  io_mmio_axi_0_w_bits_user,
  output  io_mmio_axi_0_b_ready,
  input   io_mmio_axi_0_b_valid,
  input  [1:0] io_mmio_axi_0_b_bits_resp,
  input  [4:0] io_mmio_axi_0_b_bits_id,
  input   io_mmio_axi_0_b_bits_user,
  input   io_mmio_axi_0_ar_ready,
  output  io_mmio_axi_0_ar_valid,
  output [31:0] io_mmio_axi_0_ar_bits_addr,
  output [7:0] io_mmio_axi_0_ar_bits_len,
  output [2:0] io_mmio_axi_0_ar_bits_size,
  output [1:0] io_mmio_axi_0_ar_bits_burst,
  output  io_mmio_axi_0_ar_bits_lock,
  output [3:0] io_mmio_axi_0_ar_bits_cache,
  output [2:0] io_mmio_axi_0_ar_bits_prot,
  output [3:0] io_mmio_axi_0_ar_bits_qos,
  output [3:0] io_mmio_axi_0_ar_bits_region,
  output [4:0] io_mmio_axi_0_ar_bits_id,
  output  io_mmio_axi_0_ar_bits_user,
  output  io_mmio_axi_0_r_ready,
  input   io_mmio_axi_0_r_valid,
  input  [1:0] io_mmio_axi_0_r_bits_resp,
  input  [63:0] io_mmio_axi_0_r_bits_data,
  input   io_mmio_axi_0_r_bits_last,
  input  [4:0] io_mmio_axi_0_r_bits_id,
  input   io_mmio_axi_0_r_bits_user,
  input   io_interrupts_0,
  input   io_interrupts_1,
  output  io_debugBus_req_ready,
  input   io_debugBus_req_valid,
  input  [4:0] io_debugBus_req_bits_addr,
  input  [1:0] io_debugBus_req_bits_op,
  input  [33:0] io_debugBus_req_bits_data,
  input   io_debugBus_resp_ready,
  output  io_debugBus_resp_valid,
  output [1:0] io_debugBus_resp_bits_resp,
  output [33:0] io_debugBus_resp_bits_data
);
  wire  outmemsys_clk;
  wire  outmemsys_reset;
  wire  outmemsys_io_tiles_cached_0_acquire_ready;
  wire  outmemsys_io_tiles_cached_0_acquire_valid;
  wire [25:0] outmemsys_io_tiles_cached_0_acquire_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_cached_0_acquire_bits_addr_beat;
  wire  outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_tiles_cached_0_acquire_bits_a_type;
  wire [11:0] outmemsys_io_tiles_cached_0_acquire_bits_union;
  wire [63:0] outmemsys_io_tiles_cached_0_acquire_bits_data;
  wire  outmemsys_io_tiles_cached_0_probe_ready;
  wire  outmemsys_io_tiles_cached_0_probe_valid;
  wire [25:0] outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_cached_0_probe_bits_p_type;
  wire  outmemsys_io_tiles_cached_0_release_ready;
  wire  outmemsys_io_tiles_cached_0_release_valid;
  wire [2:0] outmemsys_io_tiles_cached_0_release_bits_addr_beat;
  wire [25:0] outmemsys_io_tiles_cached_0_release_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_cached_0_release_bits_client_xact_id;
  wire  outmemsys_io_tiles_cached_0_release_bits_voluntary;
  wire [2:0] outmemsys_io_tiles_cached_0_release_bits_r_type;
  wire [63:0] outmemsys_io_tiles_cached_0_release_bits_data;
  wire  outmemsys_io_tiles_cached_0_grant_ready;
  wire  outmemsys_io_tiles_cached_0_grant_valid;
  wire [2:0] outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  wire [1:0] outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire  outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_tiles_cached_0_grant_bits_g_type;
  wire [63:0] outmemsys_io_tiles_cached_0_grant_bits_data;
  wire  outmemsys_io_tiles_cached_0_grant_bits_manager_id;
  wire  outmemsys_io_tiles_cached_0_finish_ready;
  wire  outmemsys_io_tiles_cached_0_finish_valid;
  wire [2:0] outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id;
  wire  outmemsys_io_tiles_cached_0_finish_bits_manager_id;
  wire  outmemsys_io_tiles_uncached_0_acquire_ready;
  wire  outmemsys_io_tiles_uncached_0_acquire_valid;
  wire [25:0] outmemsys_io_tiles_uncached_0_acquire_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat;
  wire  outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_tiles_uncached_0_acquire_bits_a_type;
  wire [11:0] outmemsys_io_tiles_uncached_0_acquire_bits_union;
  wire [63:0] outmemsys_io_tiles_uncached_0_acquire_bits_data;
  wire  outmemsys_io_tiles_uncached_0_grant_ready;
  wire  outmemsys_io_tiles_uncached_0_grant_valid;
  wire [2:0] outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  wire [1:0] outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire  outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  wire [63:0] outmemsys_io_tiles_uncached_0_grant_bits_data;
  wire  outmemsys_io_incoherent_0;
  wire  outmemsys_io_mem_axi_0_aw_ready;
  wire  outmemsys_io_mem_axi_0_aw_valid;
  wire [31:0] outmemsys_io_mem_axi_0_aw_bits_addr;
  wire [7:0] outmemsys_io_mem_axi_0_aw_bits_len;
  wire [2:0] outmemsys_io_mem_axi_0_aw_bits_size;
  wire [1:0] outmemsys_io_mem_axi_0_aw_bits_burst;
  wire  outmemsys_io_mem_axi_0_aw_bits_lock;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_cache;
  wire [2:0] outmemsys_io_mem_axi_0_aw_bits_prot;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_qos;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_region;
  wire [4:0] outmemsys_io_mem_axi_0_aw_bits_id;
  wire  outmemsys_io_mem_axi_0_aw_bits_user;
  wire  outmemsys_io_mem_axi_0_w_ready;
  wire  outmemsys_io_mem_axi_0_w_valid;
  wire [63:0] outmemsys_io_mem_axi_0_w_bits_data;
  wire  outmemsys_io_mem_axi_0_w_bits_last;
  wire [4:0] outmemsys_io_mem_axi_0_w_bits_id;
  wire [7:0] outmemsys_io_mem_axi_0_w_bits_strb;
  wire  outmemsys_io_mem_axi_0_w_bits_user;
  wire  outmemsys_io_mem_axi_0_b_ready;
  wire  outmemsys_io_mem_axi_0_b_valid;
  wire [1:0] outmemsys_io_mem_axi_0_b_bits_resp;
  wire [4:0] outmemsys_io_mem_axi_0_b_bits_id;
  wire  outmemsys_io_mem_axi_0_b_bits_user;
  wire  outmemsys_io_mem_axi_0_ar_ready;
  wire  outmemsys_io_mem_axi_0_ar_valid;
  wire [31:0] outmemsys_io_mem_axi_0_ar_bits_addr;
  wire [7:0] outmemsys_io_mem_axi_0_ar_bits_len;
  wire [2:0] outmemsys_io_mem_axi_0_ar_bits_size;
  wire [1:0] outmemsys_io_mem_axi_0_ar_bits_burst;
  wire  outmemsys_io_mem_axi_0_ar_bits_lock;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_cache;
  wire [2:0] outmemsys_io_mem_axi_0_ar_bits_prot;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_qos;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_region;
  wire [4:0] outmemsys_io_mem_axi_0_ar_bits_id;
  wire  outmemsys_io_mem_axi_0_ar_bits_user;
  wire  outmemsys_io_mem_axi_0_r_ready;
  wire  outmemsys_io_mem_axi_0_r_valid;
  wire [1:0] outmemsys_io_mem_axi_0_r_bits_resp;
  wire [63:0] outmemsys_io_mem_axi_0_r_bits_data;
  wire  outmemsys_io_mem_axi_0_r_bits_last;
  wire [4:0] outmemsys_io_mem_axi_0_r_bits_id;
  wire  outmemsys_io_mem_axi_0_r_bits_user;
  wire  outmemsys_io_mmio_acquire_ready;
  wire  outmemsys_io_mmio_acquire_valid;
  wire [25:0] outmemsys_io_mmio_acquire_bits_addr_block;
  wire [1:0] outmemsys_io_mmio_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_mmio_acquire_bits_addr_beat;
  wire  outmemsys_io_mmio_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_mmio_acquire_bits_a_type;
  wire [11:0] outmemsys_io_mmio_acquire_bits_union;
  wire [63:0] outmemsys_io_mmio_acquire_bits_data;
  wire  outmemsys_io_mmio_grant_ready;
  wire  outmemsys_io_mmio_grant_valid;
  wire [2:0] outmemsys_io_mmio_grant_bits_addr_beat;
  wire [1:0] outmemsys_io_mmio_grant_bits_client_xact_id;
  wire  outmemsys_io_mmio_grant_bits_manager_xact_id;
  wire  outmemsys_io_mmio_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_mmio_grant_bits_g_type;
  wire [63:0] outmemsys_io_mmio_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_clk;
  wire  TileLinkRecursiveInterconnect_2_reset;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_5_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_5_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_5_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_5_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_data;
  wire  PLIC_1_clk;
  wire  PLIC_1_reset;
  wire  PLIC_1_io_devices_0_valid;
  wire  PLIC_1_io_devices_0_ready;
  wire  PLIC_1_io_devices_0_complete;
  wire  PLIC_1_io_devices_1_valid;
  wire  PLIC_1_io_devices_1_ready;
  wire  PLIC_1_io_devices_1_complete;
  wire  PLIC_1_io_harts_0;
  wire  PLIC_1_io_harts_1;
  wire  PLIC_1_io_tl_acquire_ready;
  wire  PLIC_1_io_tl_acquire_valid;
  wire [25:0] PLIC_1_io_tl_acquire_bits_addr_block;
  wire [1:0] PLIC_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PLIC_1_io_tl_acquire_bits_addr_beat;
  wire  PLIC_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PLIC_1_io_tl_acquire_bits_a_type;
  wire [11:0] PLIC_1_io_tl_acquire_bits_union;
  wire [63:0] PLIC_1_io_tl_acquire_bits_data;
  wire  PLIC_1_io_tl_grant_ready;
  wire  PLIC_1_io_tl_grant_valid;
  wire [2:0] PLIC_1_io_tl_grant_bits_addr_beat;
  wire [1:0] PLIC_1_io_tl_grant_bits_client_xact_id;
  wire  PLIC_1_io_tl_grant_bits_manager_xact_id;
  wire  PLIC_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PLIC_1_io_tl_grant_bits_g_type;
  wire [63:0] PLIC_1_io_tl_grant_bits_data;
  wire  LevelGateway_2_clk;
  wire  LevelGateway_2_reset;
  wire  LevelGateway_2_io_interrupt;
  wire  LevelGateway_2_io_plic_valid;
  wire  LevelGateway_2_io_plic_ready;
  wire  LevelGateway_2_io_plic_complete;
  wire  LevelGateway_1_1_clk;
  wire  LevelGateway_1_1_reset;
  wire  LevelGateway_1_1_io_interrupt;
  wire  LevelGateway_1_1_io_plic_valid;
  wire  LevelGateway_1_1_io_plic_ready;
  wire  LevelGateway_1_1_io_plic_complete;
  wire  DebugModule_1_clk;
  wire  DebugModule_1_reset;
  wire  DebugModule_1_io_db_req_ready;
  wire  DebugModule_1_io_db_req_valid;
  wire [4:0] DebugModule_1_io_db_req_bits_addr;
  wire [1:0] DebugModule_1_io_db_req_bits_op;
  wire [33:0] DebugModule_1_io_db_req_bits_data;
  wire  DebugModule_1_io_db_resp_ready;
  wire  DebugModule_1_io_db_resp_valid;
  wire [1:0] DebugModule_1_io_db_resp_bits_resp;
  wire [33:0] DebugModule_1_io_db_resp_bits_data;
  wire  DebugModule_1_io_debugInterrupts_0;
  wire  DebugModule_1_io_tl_acquire_ready;
  wire  DebugModule_1_io_tl_acquire_valid;
  wire [25:0] DebugModule_1_io_tl_acquire_bits_addr_block;
  wire [1:0] DebugModule_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] DebugModule_1_io_tl_acquire_bits_addr_beat;
  wire  DebugModule_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] DebugModule_1_io_tl_acquire_bits_a_type;
  wire [11:0] DebugModule_1_io_tl_acquire_bits_union;
  wire [63:0] DebugModule_1_io_tl_acquire_bits_data;
  wire  DebugModule_1_io_tl_grant_ready;
  wire  DebugModule_1_io_tl_grant_valid;
  wire [2:0] DebugModule_1_io_tl_grant_bits_addr_beat;
  wire [1:0] DebugModule_1_io_tl_grant_bits_client_xact_id;
  wire  DebugModule_1_io_tl_grant_bits_manager_xact_id;
  wire  DebugModule_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] DebugModule_1_io_tl_grant_bits_g_type;
  wire [63:0] DebugModule_1_io_tl_grant_bits_data;
  wire  DebugModule_1_io_ndreset;
  wire  DebugModule_1_io_fullreset;
  wire  PRCI_1_clk;
  wire  PRCI_1_reset;
  wire  PRCI_1_io_interrupts_0_meip;
  wire  PRCI_1_io_interrupts_0_seip;
  wire  PRCI_1_io_interrupts_0_debug;
  wire  PRCI_1_io_tl_acquire_ready;
  wire  PRCI_1_io_tl_acquire_valid;
  wire [25:0] PRCI_1_io_tl_acquire_bits_addr_block;
  wire [1:0] PRCI_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PRCI_1_io_tl_acquire_bits_addr_beat;
  wire  PRCI_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PRCI_1_io_tl_acquire_bits_a_type;
  wire [11:0] PRCI_1_io_tl_acquire_bits_union;
  wire [63:0] PRCI_1_io_tl_acquire_bits_data;
  wire  PRCI_1_io_tl_grant_ready;
  wire  PRCI_1_io_tl_grant_valid;
  wire [2:0] PRCI_1_io_tl_grant_bits_addr_beat;
  wire [1:0] PRCI_1_io_tl_grant_bits_client_xact_id;
  wire  PRCI_1_io_tl_grant_bits_manager_xact_id;
  wire  PRCI_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PRCI_1_io_tl_grant_bits_g_type;
  wire [63:0] PRCI_1_io_tl_grant_bits_data;
  wire  PRCI_1_io_tiles_0_reset;
  wire  PRCI_1_io_tiles_0_id;
  wire  PRCI_1_io_tiles_0_interrupts_meip;
  wire  PRCI_1_io_tiles_0_interrupts_seip;
  wire  PRCI_1_io_tiles_0_interrupts_debug;
  wire  PRCI_1_io_tiles_0_interrupts_mtip;
  wire  PRCI_1_io_tiles_0_interrupts_msip;
  wire  PRCI_1_io_rtcTick;
  reg [6:0] T_8786;
  reg [31:0] GEN_2;
  wire  T_8788;
  wire [6:0] GEN_1;
  wire [7:0] T_8790;
  wire [6:0] T_8791;
  wire [6:0] GEN_0;
  wire  ROMSlave_1_clk;
  wire  ROMSlave_1_reset;
  wire  ROMSlave_1_io_acquire_ready;
  wire  ROMSlave_1_io_acquire_valid;
  wire [25:0] ROMSlave_1_io_acquire_bits_addr_block;
  wire [1:0] ROMSlave_1_io_acquire_bits_client_xact_id;
  wire [2:0] ROMSlave_1_io_acquire_bits_addr_beat;
  wire  ROMSlave_1_io_acquire_bits_is_builtin_type;
  wire [2:0] ROMSlave_1_io_acquire_bits_a_type;
  wire [11:0] ROMSlave_1_io_acquire_bits_union;
  wire [63:0] ROMSlave_1_io_acquire_bits_data;
  wire  ROMSlave_1_io_grant_ready;
  wire  ROMSlave_1_io_grant_valid;
  wire [2:0] ROMSlave_1_io_grant_bits_addr_beat;
  wire [1:0] ROMSlave_1_io_grant_bits_client_xact_id;
  wire  ROMSlave_1_io_grant_bits_manager_xact_id;
  wire  ROMSlave_1_io_grant_bits_is_builtin_type;
  wire [3:0] ROMSlave_1_io_grant_bits_g_type;
  wire [63:0] ROMSlave_1_io_grant_bits_data;
  wire  BRAMSlave_1_clk;
  wire  BRAMSlave_1_reset;
  wire  BRAMSlave_1_io_acquire_ready;
  wire  BRAMSlave_1_io_acquire_valid;
  wire [25:0] BRAMSlave_1_io_acquire_bits_addr_block;
  wire [1:0] BRAMSlave_1_io_acquire_bits_client_xact_id;
  wire [2:0] BRAMSlave_1_io_acquire_bits_addr_beat;
  wire  BRAMSlave_1_io_acquire_bits_is_builtin_type;
  wire [2:0] BRAMSlave_1_io_acquire_bits_a_type;
  wire [11:0] BRAMSlave_1_io_acquire_bits_union;
  wire [63:0] BRAMSlave_1_io_acquire_bits_data;
  wire  BRAMSlave_1_io_grant_ready;
  wire  BRAMSlave_1_io_grant_valid;
  wire [2:0] BRAMSlave_1_io_grant_bits_addr_beat;
  wire [1:0] BRAMSlave_1_io_grant_bits_client_xact_id;
  wire  BRAMSlave_1_io_grant_bits_manager_xact_id;
  wire  BRAMSlave_1_io_grant_bits_is_builtin_type;
  wire [3:0] BRAMSlave_1_io_grant_bits_g_type;
  wire [63:0] BRAMSlave_1_io_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_clk;
  wire  NastiIOTileLinkIOConverter_1_1_reset;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_acquire_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_acquire_valid;
  wire [25:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_block;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_beat;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_a_type;
  wire [11:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_union;
  wire [63:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_grant_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_grant_valid;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_addr_beat;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_client_xact_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_manager_xact_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_g_type;
  wire [63:0] NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_aw_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_aw_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_user;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_w_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_w_valid;
  wire [63:0] NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_id;
  wire [7:0] NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_strb;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_user;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_b_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_b_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_resp;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_user;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_ar_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_ar_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_user;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_r_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_r_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_resp;
  wire [63:0] NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_user;
  wire  Queue_23_1_clk;
  wire  Queue_23_1_reset;
  wire  Queue_23_1_io_enq_ready;
  wire  Queue_23_1_io_enq_valid;
  wire [31:0] Queue_23_1_io_enq_bits_addr;
  wire [7:0] Queue_23_1_io_enq_bits_len;
  wire [2:0] Queue_23_1_io_enq_bits_size;
  wire [1:0] Queue_23_1_io_enq_bits_burst;
  wire  Queue_23_1_io_enq_bits_lock;
  wire [3:0] Queue_23_1_io_enq_bits_cache;
  wire [2:0] Queue_23_1_io_enq_bits_prot;
  wire [3:0] Queue_23_1_io_enq_bits_qos;
  wire [3:0] Queue_23_1_io_enq_bits_region;
  wire [4:0] Queue_23_1_io_enq_bits_id;
  wire  Queue_23_1_io_enq_bits_user;
  wire  Queue_23_1_io_deq_ready;
  wire  Queue_23_1_io_deq_valid;
  wire [31:0] Queue_23_1_io_deq_bits_addr;
  wire [7:0] Queue_23_1_io_deq_bits_len;
  wire [2:0] Queue_23_1_io_deq_bits_size;
  wire [1:0] Queue_23_1_io_deq_bits_burst;
  wire  Queue_23_1_io_deq_bits_lock;
  wire [3:0] Queue_23_1_io_deq_bits_cache;
  wire [2:0] Queue_23_1_io_deq_bits_prot;
  wire [3:0] Queue_23_1_io_deq_bits_qos;
  wire [3:0] Queue_23_1_io_deq_bits_region;
  wire [4:0] Queue_23_1_io_deq_bits_id;
  wire  Queue_23_1_io_deq_bits_user;
  wire  Queue_23_1_io_count;
  wire  Queue_24_1_clk;
  wire  Queue_24_1_reset;
  wire  Queue_24_1_io_enq_ready;
  wire  Queue_24_1_io_enq_valid;
  wire [31:0] Queue_24_1_io_enq_bits_addr;
  wire [7:0] Queue_24_1_io_enq_bits_len;
  wire [2:0] Queue_24_1_io_enq_bits_size;
  wire [1:0] Queue_24_1_io_enq_bits_burst;
  wire  Queue_24_1_io_enq_bits_lock;
  wire [3:0] Queue_24_1_io_enq_bits_cache;
  wire [2:0] Queue_24_1_io_enq_bits_prot;
  wire [3:0] Queue_24_1_io_enq_bits_qos;
  wire [3:0] Queue_24_1_io_enq_bits_region;
  wire [4:0] Queue_24_1_io_enq_bits_id;
  wire  Queue_24_1_io_enq_bits_user;
  wire  Queue_24_1_io_deq_ready;
  wire  Queue_24_1_io_deq_valid;
  wire [31:0] Queue_24_1_io_deq_bits_addr;
  wire [7:0] Queue_24_1_io_deq_bits_len;
  wire [2:0] Queue_24_1_io_deq_bits_size;
  wire [1:0] Queue_24_1_io_deq_bits_burst;
  wire  Queue_24_1_io_deq_bits_lock;
  wire [3:0] Queue_24_1_io_deq_bits_cache;
  wire [2:0] Queue_24_1_io_deq_bits_prot;
  wire [3:0] Queue_24_1_io_deq_bits_qos;
  wire [3:0] Queue_24_1_io_deq_bits_region;
  wire [4:0] Queue_24_1_io_deq_bits_id;
  wire  Queue_24_1_io_deq_bits_user;
  wire  Queue_24_1_io_count;
  wire  Queue_25_1_clk;
  wire  Queue_25_1_reset;
  wire  Queue_25_1_io_enq_ready;
  wire  Queue_25_1_io_enq_valid;
  wire [63:0] Queue_25_1_io_enq_bits_data;
  wire  Queue_25_1_io_enq_bits_last;
  wire [4:0] Queue_25_1_io_enq_bits_id;
  wire [7:0] Queue_25_1_io_enq_bits_strb;
  wire  Queue_25_1_io_enq_bits_user;
  wire  Queue_25_1_io_deq_ready;
  wire  Queue_25_1_io_deq_valid;
  wire [63:0] Queue_25_1_io_deq_bits_data;
  wire  Queue_25_1_io_deq_bits_last;
  wire [4:0] Queue_25_1_io_deq_bits_id;
  wire [7:0] Queue_25_1_io_deq_bits_strb;
  wire  Queue_25_1_io_deq_bits_user;
  wire [1:0] Queue_25_1_io_count;
  wire  Queue_26_1_clk;
  wire  Queue_26_1_reset;
  wire  Queue_26_1_io_enq_ready;
  wire  Queue_26_1_io_enq_valid;
  wire [1:0] Queue_26_1_io_enq_bits_resp;
  wire [63:0] Queue_26_1_io_enq_bits_data;
  wire  Queue_26_1_io_enq_bits_last;
  wire [4:0] Queue_26_1_io_enq_bits_id;
  wire  Queue_26_1_io_enq_bits_user;
  wire  Queue_26_1_io_deq_ready;
  wire  Queue_26_1_io_deq_valid;
  wire [1:0] Queue_26_1_io_deq_bits_resp;
  wire [63:0] Queue_26_1_io_deq_bits_data;
  wire  Queue_26_1_io_deq_bits_last;
  wire [4:0] Queue_26_1_io_deq_bits_id;
  wire  Queue_26_1_io_deq_bits_user;
  wire [1:0] Queue_26_1_io_count;
  wire  Queue_27_1_clk;
  wire  Queue_27_1_reset;
  wire  Queue_27_1_io_enq_ready;
  wire  Queue_27_1_io_enq_valid;
  wire [1:0] Queue_27_1_io_enq_bits_resp;
  wire [4:0] Queue_27_1_io_enq_bits_id;
  wire  Queue_27_1_io_enq_bits_user;
  wire  Queue_27_1_io_deq_ready;
  wire  Queue_27_1_io_deq_valid;
  wire [1:0] Queue_27_1_io_deq_bits_resp;
  wire [4:0] Queue_27_1_io_deq_bits_id;
  wire  Queue_27_1_io_deq_bits_user;
  wire  Queue_27_1_io_count;
  OuterMemorySystem outmemsys (
    .clk(outmemsys_clk),
    .reset(outmemsys_reset),
    .io_tiles_cached_0_acquire_ready(outmemsys_io_tiles_cached_0_acquire_ready),
    .io_tiles_cached_0_acquire_valid(outmemsys_io_tiles_cached_0_acquire_valid),
    .io_tiles_cached_0_acquire_bits_addr_block(outmemsys_io_tiles_cached_0_acquire_bits_addr_block),
    .io_tiles_cached_0_acquire_bits_client_xact_id(outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id),
    .io_tiles_cached_0_acquire_bits_addr_beat(outmemsys_io_tiles_cached_0_acquire_bits_addr_beat),
    .io_tiles_cached_0_acquire_bits_is_builtin_type(outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type),
    .io_tiles_cached_0_acquire_bits_a_type(outmemsys_io_tiles_cached_0_acquire_bits_a_type),
    .io_tiles_cached_0_acquire_bits_union(outmemsys_io_tiles_cached_0_acquire_bits_union),
    .io_tiles_cached_0_acquire_bits_data(outmemsys_io_tiles_cached_0_acquire_bits_data),
    .io_tiles_cached_0_probe_ready(outmemsys_io_tiles_cached_0_probe_ready),
    .io_tiles_cached_0_probe_valid(outmemsys_io_tiles_cached_0_probe_valid),
    .io_tiles_cached_0_probe_bits_addr_block(outmemsys_io_tiles_cached_0_probe_bits_addr_block),
    .io_tiles_cached_0_probe_bits_p_type(outmemsys_io_tiles_cached_0_probe_bits_p_type),
    .io_tiles_cached_0_release_ready(outmemsys_io_tiles_cached_0_release_ready),
    .io_tiles_cached_0_release_valid(outmemsys_io_tiles_cached_0_release_valid),
    .io_tiles_cached_0_release_bits_addr_beat(outmemsys_io_tiles_cached_0_release_bits_addr_beat),
    .io_tiles_cached_0_release_bits_addr_block(outmemsys_io_tiles_cached_0_release_bits_addr_block),
    .io_tiles_cached_0_release_bits_client_xact_id(outmemsys_io_tiles_cached_0_release_bits_client_xact_id),
    .io_tiles_cached_0_release_bits_voluntary(outmemsys_io_tiles_cached_0_release_bits_voluntary),
    .io_tiles_cached_0_release_bits_r_type(outmemsys_io_tiles_cached_0_release_bits_r_type),
    .io_tiles_cached_0_release_bits_data(outmemsys_io_tiles_cached_0_release_bits_data),
    .io_tiles_cached_0_grant_ready(outmemsys_io_tiles_cached_0_grant_ready),
    .io_tiles_cached_0_grant_valid(outmemsys_io_tiles_cached_0_grant_valid),
    .io_tiles_cached_0_grant_bits_addr_beat(outmemsys_io_tiles_cached_0_grant_bits_addr_beat),
    .io_tiles_cached_0_grant_bits_client_xact_id(outmemsys_io_tiles_cached_0_grant_bits_client_xact_id),
    .io_tiles_cached_0_grant_bits_manager_xact_id(outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id),
    .io_tiles_cached_0_grant_bits_is_builtin_type(outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type),
    .io_tiles_cached_0_grant_bits_g_type(outmemsys_io_tiles_cached_0_grant_bits_g_type),
    .io_tiles_cached_0_grant_bits_data(outmemsys_io_tiles_cached_0_grant_bits_data),
    .io_tiles_cached_0_grant_bits_manager_id(outmemsys_io_tiles_cached_0_grant_bits_manager_id),
    .io_tiles_cached_0_finish_ready(outmemsys_io_tiles_cached_0_finish_ready),
    .io_tiles_cached_0_finish_valid(outmemsys_io_tiles_cached_0_finish_valid),
    .io_tiles_cached_0_finish_bits_manager_xact_id(outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id),
    .io_tiles_cached_0_finish_bits_manager_id(outmemsys_io_tiles_cached_0_finish_bits_manager_id),
    .io_tiles_uncached_0_acquire_ready(outmemsys_io_tiles_uncached_0_acquire_ready),
    .io_tiles_uncached_0_acquire_valid(outmemsys_io_tiles_uncached_0_acquire_valid),
    .io_tiles_uncached_0_acquire_bits_addr_block(outmemsys_io_tiles_uncached_0_acquire_bits_addr_block),
    .io_tiles_uncached_0_acquire_bits_client_xact_id(outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id),
    .io_tiles_uncached_0_acquire_bits_addr_beat(outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat),
    .io_tiles_uncached_0_acquire_bits_is_builtin_type(outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type),
    .io_tiles_uncached_0_acquire_bits_a_type(outmemsys_io_tiles_uncached_0_acquire_bits_a_type),
    .io_tiles_uncached_0_acquire_bits_union(outmemsys_io_tiles_uncached_0_acquire_bits_union),
    .io_tiles_uncached_0_acquire_bits_data(outmemsys_io_tiles_uncached_0_acquire_bits_data),
    .io_tiles_uncached_0_grant_ready(outmemsys_io_tiles_uncached_0_grant_ready),
    .io_tiles_uncached_0_grant_valid(outmemsys_io_tiles_uncached_0_grant_valid),
    .io_tiles_uncached_0_grant_bits_addr_beat(outmemsys_io_tiles_uncached_0_grant_bits_addr_beat),
    .io_tiles_uncached_0_grant_bits_client_xact_id(outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id),
    .io_tiles_uncached_0_grant_bits_manager_xact_id(outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id),
    .io_tiles_uncached_0_grant_bits_is_builtin_type(outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type),
    .io_tiles_uncached_0_grant_bits_g_type(outmemsys_io_tiles_uncached_0_grant_bits_g_type),
    .io_tiles_uncached_0_grant_bits_data(outmemsys_io_tiles_uncached_0_grant_bits_data),
    .io_incoherent_0(outmemsys_io_incoherent_0),
    .io_mem_axi_0_aw_ready(outmemsys_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(outmemsys_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(outmemsys_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(outmemsys_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(outmemsys_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(outmemsys_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(outmemsys_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(outmemsys_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(outmemsys_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(outmemsys_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(outmemsys_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(outmemsys_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(outmemsys_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(outmemsys_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(outmemsys_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(outmemsys_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(outmemsys_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(outmemsys_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(outmemsys_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(outmemsys_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(outmemsys_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(outmemsys_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(outmemsys_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(outmemsys_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(outmemsys_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(outmemsys_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(outmemsys_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(outmemsys_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(outmemsys_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(outmemsys_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(outmemsys_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(outmemsys_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(outmemsys_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(outmemsys_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(outmemsys_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(outmemsys_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(outmemsys_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(outmemsys_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(outmemsys_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(outmemsys_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(outmemsys_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(outmemsys_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(outmemsys_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(outmemsys_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(outmemsys_io_mem_axi_0_r_bits_user),
    .io_mmio_acquire_ready(outmemsys_io_mmio_acquire_ready),
    .io_mmio_acquire_valid(outmemsys_io_mmio_acquire_valid),
    .io_mmio_acquire_bits_addr_block(outmemsys_io_mmio_acquire_bits_addr_block),
    .io_mmio_acquire_bits_client_xact_id(outmemsys_io_mmio_acquire_bits_client_xact_id),
    .io_mmio_acquire_bits_addr_beat(outmemsys_io_mmio_acquire_bits_addr_beat),
    .io_mmio_acquire_bits_is_builtin_type(outmemsys_io_mmio_acquire_bits_is_builtin_type),
    .io_mmio_acquire_bits_a_type(outmemsys_io_mmio_acquire_bits_a_type),
    .io_mmio_acquire_bits_union(outmemsys_io_mmio_acquire_bits_union),
    .io_mmio_acquire_bits_data(outmemsys_io_mmio_acquire_bits_data),
    .io_mmio_grant_ready(outmemsys_io_mmio_grant_ready),
    .io_mmio_grant_valid(outmemsys_io_mmio_grant_valid),
    .io_mmio_grant_bits_addr_beat(outmemsys_io_mmio_grant_bits_addr_beat),
    .io_mmio_grant_bits_client_xact_id(outmemsys_io_mmio_grant_bits_client_xact_id),
    .io_mmio_grant_bits_manager_xact_id(outmemsys_io_mmio_grant_bits_manager_xact_id),
    .io_mmio_grant_bits_is_builtin_type(outmemsys_io_mmio_grant_bits_is_builtin_type),
    .io_mmio_grant_bits_g_type(outmemsys_io_mmio_grant_bits_g_type),
    .io_mmio_grant_bits_data(outmemsys_io_mmio_grant_bits_data)
  );
  TileLinkRecursiveInterconnect TileLinkRecursiveInterconnect_2 (
    .clk(TileLinkRecursiveInterconnect_2_clk),
    .reset(TileLinkRecursiveInterconnect_2_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_2_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_2_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_2_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_2_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_2_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_2_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_2_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_2_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_2_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_2_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(TileLinkRecursiveInterconnect_2_io_out_4_grant_ready),
    .io_out_4_grant_valid(TileLinkRecursiveInterconnect_2_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_data),
    .io_out_5_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_5_acquire_ready),
    .io_out_5_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_5_acquire_valid),
    .io_out_5_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_addr_block),
    .io_out_5_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_client_xact_id),
    .io_out_5_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_addr_beat),
    .io_out_5_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_is_builtin_type),
    .io_out_5_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_a_type),
    .io_out_5_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_union),
    .io_out_5_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_data),
    .io_out_5_grant_ready(TileLinkRecursiveInterconnect_2_io_out_5_grant_ready),
    .io_out_5_grant_valid(TileLinkRecursiveInterconnect_2_io_out_5_grant_valid),
    .io_out_5_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_addr_beat),
    .io_out_5_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_client_xact_id),
    .io_out_5_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_manager_xact_id),
    .io_out_5_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_is_builtin_type),
    .io_out_5_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_g_type),
    .io_out_5_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_data)
  );
  PLIC PLIC_1 (
    .clk(PLIC_1_clk),
    .reset(PLIC_1_reset),
    .io_devices_0_valid(PLIC_1_io_devices_0_valid),
    .io_devices_0_ready(PLIC_1_io_devices_0_ready),
    .io_devices_0_complete(PLIC_1_io_devices_0_complete),
    .io_devices_1_valid(PLIC_1_io_devices_1_valid),
    .io_devices_1_ready(PLIC_1_io_devices_1_ready),
    .io_devices_1_complete(PLIC_1_io_devices_1_complete),
    .io_harts_0(PLIC_1_io_harts_0),
    .io_harts_1(PLIC_1_io_harts_1),
    .io_tl_acquire_ready(PLIC_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(PLIC_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PLIC_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PLIC_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PLIC_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PLIC_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PLIC_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PLIC_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PLIC_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PLIC_1_io_tl_grant_ready),
    .io_tl_grant_valid(PLIC_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PLIC_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PLIC_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PLIC_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PLIC_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PLIC_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PLIC_1_io_tl_grant_bits_data)
  );
  LevelGateway LevelGateway_2 (
    .clk(LevelGateway_2_clk),
    .reset(LevelGateway_2_reset),
    .io_interrupt(LevelGateway_2_io_interrupt),
    .io_plic_valid(LevelGateway_2_io_plic_valid),
    .io_plic_ready(LevelGateway_2_io_plic_ready),
    .io_plic_complete(LevelGateway_2_io_plic_complete)
  );
  LevelGateway LevelGateway_1_1 (
    .clk(LevelGateway_1_1_clk),
    .reset(LevelGateway_1_1_reset),
    .io_interrupt(LevelGateway_1_1_io_interrupt),
    .io_plic_valid(LevelGateway_1_1_io_plic_valid),
    .io_plic_ready(LevelGateway_1_1_io_plic_ready),
    .io_plic_complete(LevelGateway_1_1_io_plic_complete)
  );
  DebugModule DebugModule_1 (
    .clk(DebugModule_1_clk),
    .reset(DebugModule_1_reset),
    .io_db_req_ready(DebugModule_1_io_db_req_ready),
    .io_db_req_valid(DebugModule_1_io_db_req_valid),
    .io_db_req_bits_addr(DebugModule_1_io_db_req_bits_addr),
    .io_db_req_bits_op(DebugModule_1_io_db_req_bits_op),
    .io_db_req_bits_data(DebugModule_1_io_db_req_bits_data),
    .io_db_resp_ready(DebugModule_1_io_db_resp_ready),
    .io_db_resp_valid(DebugModule_1_io_db_resp_valid),
    .io_db_resp_bits_resp(DebugModule_1_io_db_resp_bits_resp),
    .io_db_resp_bits_data(DebugModule_1_io_db_resp_bits_data),
    .io_debugInterrupts_0(DebugModule_1_io_debugInterrupts_0),
    .io_tl_acquire_ready(DebugModule_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(DebugModule_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(DebugModule_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(DebugModule_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(DebugModule_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(DebugModule_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(DebugModule_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(DebugModule_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(DebugModule_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(DebugModule_1_io_tl_grant_ready),
    .io_tl_grant_valid(DebugModule_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(DebugModule_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(DebugModule_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(DebugModule_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(DebugModule_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(DebugModule_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(DebugModule_1_io_tl_grant_bits_data),
    .io_ndreset(DebugModule_1_io_ndreset),
    .io_fullreset(DebugModule_1_io_fullreset)
  );
  PRCI PRCI_1 (
    .clk(PRCI_1_clk),
    .reset(PRCI_1_reset),
    .io_interrupts_0_meip(PRCI_1_io_interrupts_0_meip),
    .io_interrupts_0_seip(PRCI_1_io_interrupts_0_seip),
    .io_interrupts_0_debug(PRCI_1_io_interrupts_0_debug),
    .io_tl_acquire_ready(PRCI_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(PRCI_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PRCI_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PRCI_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PRCI_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PRCI_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PRCI_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PRCI_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PRCI_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PRCI_1_io_tl_grant_ready),
    .io_tl_grant_valid(PRCI_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PRCI_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PRCI_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PRCI_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PRCI_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PRCI_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PRCI_1_io_tl_grant_bits_data),
    .io_tiles_0_reset(PRCI_1_io_tiles_0_reset),
    .io_tiles_0_id(PRCI_1_io_tiles_0_id),
    .io_tiles_0_interrupts_meip(PRCI_1_io_tiles_0_interrupts_meip),
    .io_tiles_0_interrupts_seip(PRCI_1_io_tiles_0_interrupts_seip),
    .io_tiles_0_interrupts_debug(PRCI_1_io_tiles_0_interrupts_debug),
    .io_tiles_0_interrupts_mtip(PRCI_1_io_tiles_0_interrupts_mtip),
    .io_tiles_0_interrupts_msip(PRCI_1_io_tiles_0_interrupts_msip),
    .io_rtcTick(PRCI_1_io_rtcTick)
  );
  ROMSlave ROMSlave_1 (
    .clk(ROMSlave_1_clk),
    .reset(ROMSlave_1_reset),
    .io_acquire_ready(ROMSlave_1_io_acquire_ready),
    .io_acquire_valid(ROMSlave_1_io_acquire_valid),
    .io_acquire_bits_addr_block(ROMSlave_1_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(ROMSlave_1_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(ROMSlave_1_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(ROMSlave_1_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(ROMSlave_1_io_acquire_bits_a_type),
    .io_acquire_bits_union(ROMSlave_1_io_acquire_bits_union),
    .io_acquire_bits_data(ROMSlave_1_io_acquire_bits_data),
    .io_grant_ready(ROMSlave_1_io_grant_ready),
    .io_grant_valid(ROMSlave_1_io_grant_valid),
    .io_grant_bits_addr_beat(ROMSlave_1_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(ROMSlave_1_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(ROMSlave_1_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(ROMSlave_1_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(ROMSlave_1_io_grant_bits_g_type),
    .io_grant_bits_data(ROMSlave_1_io_grant_bits_data)
  );
  BRAMSlave BRAMSlave_1 (
    .clk(BRAMSlave_1_clk),
    .reset(BRAMSlave_1_reset),
    .io_acquire_ready(BRAMSlave_1_io_acquire_ready),
    .io_acquire_valid(BRAMSlave_1_io_acquire_valid),
    .io_acquire_bits_addr_block(BRAMSlave_1_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(BRAMSlave_1_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(BRAMSlave_1_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(BRAMSlave_1_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(BRAMSlave_1_io_acquire_bits_a_type),
    .io_acquire_bits_union(BRAMSlave_1_io_acquire_bits_union),
    .io_acquire_bits_data(BRAMSlave_1_io_acquire_bits_data),
    .io_grant_ready(BRAMSlave_1_io_grant_ready),
    .io_grant_valid(BRAMSlave_1_io_grant_valid),
    .io_grant_bits_addr_beat(BRAMSlave_1_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(BRAMSlave_1_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(BRAMSlave_1_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(BRAMSlave_1_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(BRAMSlave_1_io_grant_bits_g_type),
    .io_grant_bits_data(BRAMSlave_1_io_grant_bits_data)
  );
  NastiIOTileLinkIOConverter_1 NastiIOTileLinkIOConverter_1_1 (
    .clk(NastiIOTileLinkIOConverter_1_1_clk),
    .reset(NastiIOTileLinkIOConverter_1_1_reset),
    .io_tl_acquire_ready(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(NastiIOTileLinkIOConverter_1_1_io_tl_grant_ready),
    .io_tl_grant_valid(NastiIOTileLinkIOConverter_1_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_data),
    .io_nasti_aw_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_ready),
    .io_nasti_aw_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_user),
    .io_nasti_w_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_w_ready),
    .io_nasti_w_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_w_valid),
    .io_nasti_w_bits_data(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_user),
    .io_nasti_b_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_b_ready),
    .io_nasti_b_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_b_valid),
    .io_nasti_b_bits_resp(NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_user),
    .io_nasti_ar_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_ready),
    .io_nasti_ar_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_user),
    .io_nasti_r_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_r_ready),
    .io_nasti_r_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_r_valid),
    .io_nasti_r_bits_resp(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_user)
  );
  Queue_15 Queue_23_1 (
    .clk(Queue_23_1_clk),
    .reset(Queue_23_1_reset),
    .io_enq_ready(Queue_23_1_io_enq_ready),
    .io_enq_valid(Queue_23_1_io_enq_valid),
    .io_enq_bits_addr(Queue_23_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_23_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_23_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_23_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_23_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_23_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_23_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_23_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_23_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_23_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_23_1_io_enq_bits_user),
    .io_deq_ready(Queue_23_1_io_deq_ready),
    .io_deq_valid(Queue_23_1_io_deq_valid),
    .io_deq_bits_addr(Queue_23_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_23_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_23_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_23_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_23_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_23_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_23_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_23_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_23_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_23_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_23_1_io_deq_bits_user),
    .io_count(Queue_23_1_io_count)
  );
  Queue_15 Queue_24_1 (
    .clk(Queue_24_1_clk),
    .reset(Queue_24_1_reset),
    .io_enq_ready(Queue_24_1_io_enq_ready),
    .io_enq_valid(Queue_24_1_io_enq_valid),
    .io_enq_bits_addr(Queue_24_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_24_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_24_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_24_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_24_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_24_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_24_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_24_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_24_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_24_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_24_1_io_enq_bits_user),
    .io_deq_ready(Queue_24_1_io_deq_ready),
    .io_deq_valid(Queue_24_1_io_deq_valid),
    .io_deq_bits_addr(Queue_24_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_24_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_24_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_24_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_24_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_24_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_24_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_24_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_24_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_24_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_24_1_io_deq_bits_user),
    .io_count(Queue_24_1_io_count)
  );
  Queue_17 Queue_25_1 (
    .clk(Queue_25_1_clk),
    .reset(Queue_25_1_reset),
    .io_enq_ready(Queue_25_1_io_enq_ready),
    .io_enq_valid(Queue_25_1_io_enq_valid),
    .io_enq_bits_data(Queue_25_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_25_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_25_1_io_enq_bits_id),
    .io_enq_bits_strb(Queue_25_1_io_enq_bits_strb),
    .io_enq_bits_user(Queue_25_1_io_enq_bits_user),
    .io_deq_ready(Queue_25_1_io_deq_ready),
    .io_deq_valid(Queue_25_1_io_deq_valid),
    .io_deq_bits_data(Queue_25_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_25_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_25_1_io_deq_bits_id),
    .io_deq_bits_strb(Queue_25_1_io_deq_bits_strb),
    .io_deq_bits_user(Queue_25_1_io_deq_bits_user),
    .io_count(Queue_25_1_io_count)
  );
  Queue_18 Queue_26_1 (
    .clk(Queue_26_1_clk),
    .reset(Queue_26_1_reset),
    .io_enq_ready(Queue_26_1_io_enq_ready),
    .io_enq_valid(Queue_26_1_io_enq_valid),
    .io_enq_bits_resp(Queue_26_1_io_enq_bits_resp),
    .io_enq_bits_data(Queue_26_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_26_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_26_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_26_1_io_enq_bits_user),
    .io_deq_ready(Queue_26_1_io_deq_ready),
    .io_deq_valid(Queue_26_1_io_deq_valid),
    .io_deq_bits_resp(Queue_26_1_io_deq_bits_resp),
    .io_deq_bits_data(Queue_26_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_26_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_26_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_26_1_io_deq_bits_user),
    .io_count(Queue_26_1_io_count)
  );
  Queue_19 Queue_27_1 (
    .clk(Queue_27_1_clk),
    .reset(Queue_27_1_reset),
    .io_enq_ready(Queue_27_1_io_enq_ready),
    .io_enq_valid(Queue_27_1_io_enq_valid),
    .io_enq_bits_resp(Queue_27_1_io_enq_bits_resp),
    .io_enq_bits_id(Queue_27_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_27_1_io_enq_bits_user),
    .io_deq_ready(Queue_27_1_io_deq_ready),
    .io_deq_valid(Queue_27_1_io_deq_valid),
    .io_deq_bits_resp(Queue_27_1_io_deq_bits_resp),
    .io_deq_bits_id(Queue_27_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_27_1_io_deq_bits_user),
    .io_count(Queue_27_1_io_count)
  );
  assign io_mem_axi_0_aw_valid = outmemsys_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = outmemsys_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = outmemsys_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = outmemsys_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = outmemsys_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = outmemsys_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = outmemsys_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = outmemsys_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = outmemsys_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = outmemsys_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = outmemsys_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = outmemsys_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = outmemsys_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = outmemsys_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = outmemsys_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = outmemsys_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = outmemsys_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = outmemsys_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = outmemsys_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = outmemsys_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = outmemsys_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = outmemsys_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = outmemsys_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = outmemsys_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = outmemsys_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = outmemsys_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = outmemsys_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = outmemsys_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = outmemsys_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = outmemsys_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = outmemsys_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = outmemsys_io_mem_axi_0_r_ready;
  assign io_tiles_cached_0_acquire_ready = outmemsys_io_tiles_cached_0_acquire_ready;
  assign io_tiles_cached_0_probe_valid = outmemsys_io_tiles_cached_0_probe_valid;
  assign io_tiles_cached_0_probe_bits_addr_block = outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_bits_p_type = outmemsys_io_tiles_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_release_ready = outmemsys_io_tiles_cached_0_release_ready;
  assign io_tiles_cached_0_grant_valid = outmemsys_io_tiles_cached_0_grant_valid;
  assign io_tiles_cached_0_grant_bits_addr_beat = outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_bits_client_xact_id = outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_g_type = outmemsys_io_tiles_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_data = outmemsys_io_tiles_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_manager_id = outmemsys_io_tiles_cached_0_grant_bits_manager_id;
  assign io_tiles_cached_0_finish_ready = outmemsys_io_tiles_cached_0_finish_ready;
  assign io_tiles_uncached_0_acquire_ready = outmemsys_io_tiles_uncached_0_acquire_ready;
  assign io_tiles_uncached_0_grant_valid = outmemsys_io_tiles_uncached_0_grant_valid;
  assign io_tiles_uncached_0_grant_bits_addr_beat = outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_g_type = outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_data = outmemsys_io_tiles_uncached_0_grant_bits_data;
  assign io_prci_0_reset = reset;
  assign io_prci_0_id = PRCI_1_io_tiles_0_id;
  assign io_prci_0_interrupts_meip = PRCI_1_io_tiles_0_interrupts_meip;
  assign io_prci_0_interrupts_seip = PRCI_1_io_tiles_0_interrupts_seip;
  assign io_prci_0_interrupts_debug = PRCI_1_io_tiles_0_interrupts_debug;
  assign io_prci_0_interrupts_mtip = PRCI_1_io_tiles_0_interrupts_mtip;
  assign io_prci_0_interrupts_msip = PRCI_1_io_tiles_0_interrupts_msip;
  assign io_mmio_axi_0_aw_valid = Queue_24_1_io_deq_valid;
  assign io_mmio_axi_0_aw_bits_addr = Queue_24_1_io_deq_bits_addr;
  assign io_mmio_axi_0_aw_bits_len = Queue_24_1_io_deq_bits_len;
  assign io_mmio_axi_0_aw_bits_size = Queue_24_1_io_deq_bits_size;
  assign io_mmio_axi_0_aw_bits_burst = Queue_24_1_io_deq_bits_burst;
  assign io_mmio_axi_0_aw_bits_lock = Queue_24_1_io_deq_bits_lock;
  assign io_mmio_axi_0_aw_bits_cache = Queue_24_1_io_deq_bits_cache;
  assign io_mmio_axi_0_aw_bits_prot = Queue_24_1_io_deq_bits_prot;
  assign io_mmio_axi_0_aw_bits_qos = Queue_24_1_io_deq_bits_qos;
  assign io_mmio_axi_0_aw_bits_region = Queue_24_1_io_deq_bits_region;
  assign io_mmio_axi_0_aw_bits_id = Queue_24_1_io_deq_bits_id;
  assign io_mmio_axi_0_aw_bits_user = Queue_24_1_io_deq_bits_user;
  assign io_mmio_axi_0_w_valid = Queue_25_1_io_deq_valid;
  assign io_mmio_axi_0_w_bits_data = Queue_25_1_io_deq_bits_data;
  assign io_mmio_axi_0_w_bits_last = Queue_25_1_io_deq_bits_last;
  assign io_mmio_axi_0_w_bits_id = Queue_25_1_io_deq_bits_id;
  assign io_mmio_axi_0_w_bits_strb = Queue_25_1_io_deq_bits_strb;
  assign io_mmio_axi_0_w_bits_user = Queue_25_1_io_deq_bits_user;
  assign io_mmio_axi_0_b_ready = Queue_27_1_io_enq_ready;
  assign io_mmio_axi_0_ar_valid = Queue_23_1_io_deq_valid;
  assign io_mmio_axi_0_ar_bits_addr = Queue_23_1_io_deq_bits_addr;
  assign io_mmio_axi_0_ar_bits_len = Queue_23_1_io_deq_bits_len;
  assign io_mmio_axi_0_ar_bits_size = Queue_23_1_io_deq_bits_size;
  assign io_mmio_axi_0_ar_bits_burst = Queue_23_1_io_deq_bits_burst;
  assign io_mmio_axi_0_ar_bits_lock = Queue_23_1_io_deq_bits_lock;
  assign io_mmio_axi_0_ar_bits_cache = Queue_23_1_io_deq_bits_cache;
  assign io_mmio_axi_0_ar_bits_prot = Queue_23_1_io_deq_bits_prot;
  assign io_mmio_axi_0_ar_bits_qos = Queue_23_1_io_deq_bits_qos;
  assign io_mmio_axi_0_ar_bits_region = Queue_23_1_io_deq_bits_region;
  assign io_mmio_axi_0_ar_bits_id = Queue_23_1_io_deq_bits_id;
  assign io_mmio_axi_0_ar_bits_user = Queue_23_1_io_deq_bits_user;
  assign io_mmio_axi_0_r_ready = Queue_26_1_io_enq_ready;
  assign io_debugBus_req_ready = DebugModule_1_io_db_req_ready;
  assign io_debugBus_resp_valid = DebugModule_1_io_db_resp_valid;
  assign io_debugBus_resp_bits_resp = DebugModule_1_io_db_resp_bits_resp;
  assign io_debugBus_resp_bits_data = DebugModule_1_io_db_resp_bits_data;
  assign outmemsys_clk = clk;
  assign outmemsys_reset = reset;
  assign outmemsys_io_tiles_cached_0_acquire_valid = io_tiles_cached_0_acquire_valid;
  assign outmemsys_io_tiles_cached_0_acquire_bits_addr_block = io_tiles_cached_0_acquire_bits_addr_block;
  assign outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id = io_tiles_cached_0_acquire_bits_client_xact_id;
  assign outmemsys_io_tiles_cached_0_acquire_bits_addr_beat = io_tiles_cached_0_acquire_bits_addr_beat;
  assign outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type = io_tiles_cached_0_acquire_bits_is_builtin_type;
  assign outmemsys_io_tiles_cached_0_acquire_bits_a_type = io_tiles_cached_0_acquire_bits_a_type;
  assign outmemsys_io_tiles_cached_0_acquire_bits_union = io_tiles_cached_0_acquire_bits_union;
  assign outmemsys_io_tiles_cached_0_acquire_bits_data = io_tiles_cached_0_acquire_bits_data;
  assign outmemsys_io_tiles_cached_0_probe_ready = io_tiles_cached_0_probe_ready;
  assign outmemsys_io_tiles_cached_0_release_valid = io_tiles_cached_0_release_valid;
  assign outmemsys_io_tiles_cached_0_release_bits_addr_beat = io_tiles_cached_0_release_bits_addr_beat;
  assign outmemsys_io_tiles_cached_0_release_bits_addr_block = io_tiles_cached_0_release_bits_addr_block;
  assign outmemsys_io_tiles_cached_0_release_bits_client_xact_id = io_tiles_cached_0_release_bits_client_xact_id;
  assign outmemsys_io_tiles_cached_0_release_bits_voluntary = io_tiles_cached_0_release_bits_voluntary;
  assign outmemsys_io_tiles_cached_0_release_bits_r_type = io_tiles_cached_0_release_bits_r_type;
  assign outmemsys_io_tiles_cached_0_release_bits_data = io_tiles_cached_0_release_bits_data;
  assign outmemsys_io_tiles_cached_0_grant_ready = io_tiles_cached_0_grant_ready;
  assign outmemsys_io_tiles_cached_0_finish_valid = io_tiles_cached_0_finish_valid;
  assign outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id = io_tiles_cached_0_finish_bits_manager_xact_id;
  assign outmemsys_io_tiles_cached_0_finish_bits_manager_id = io_tiles_cached_0_finish_bits_manager_id;
  assign outmemsys_io_tiles_uncached_0_acquire_valid = io_tiles_uncached_0_acquire_valid;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_addr_block = io_tiles_uncached_0_acquire_bits_addr_block;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id = io_tiles_uncached_0_acquire_bits_client_xact_id;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat = io_tiles_uncached_0_acquire_bits_addr_beat;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type = io_tiles_uncached_0_acquire_bits_is_builtin_type;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_a_type = io_tiles_uncached_0_acquire_bits_a_type;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_union = io_tiles_uncached_0_acquire_bits_union;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_data = io_tiles_uncached_0_acquire_bits_data;
  assign outmemsys_io_tiles_uncached_0_grant_ready = io_tiles_uncached_0_grant_ready;
  assign outmemsys_io_incoherent_0 = 1'h0;
  assign outmemsys_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign outmemsys_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign outmemsys_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign outmemsys_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign outmemsys_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign outmemsys_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign outmemsys_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign outmemsys_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign outmemsys_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign outmemsys_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign outmemsys_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign outmemsys_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign outmemsys_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign outmemsys_io_mmio_acquire_ready = TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready;
  assign outmemsys_io_mmio_grant_valid = TileLinkRecursiveInterconnect_2_io_in_0_grant_valid;
  assign outmemsys_io_mmio_grant_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat;
  assign outmemsys_io_mmio_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id;
  assign outmemsys_io_mmio_grant_bits_manager_xact_id = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id;
  assign outmemsys_io_mmio_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type;
  assign outmemsys_io_mmio_grant_bits_g_type = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type;
  assign outmemsys_io_mmio_grant_bits_data = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_clk = clk;
  assign TileLinkRecursiveInterconnect_2_reset = reset;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid = outmemsys_io_mmio_acquire_valid;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block = outmemsys_io_mmio_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id = outmemsys_io_mmio_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat = outmemsys_io_mmio_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type = outmemsys_io_mmio_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type = outmemsys_io_mmio_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union = outmemsys_io_mmio_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data = outmemsys_io_mmio_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_in_0_grant_ready = outmemsys_io_mmio_grant_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready = DebugModule_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_valid = DebugModule_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat = DebugModule_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id = DebugModule_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id = DebugModule_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type = DebugModule_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type = DebugModule_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data = DebugModule_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready = ROMSlave_1_io_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_valid = ROMSlave_1_io_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat = ROMSlave_1_io_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id = ROMSlave_1_io_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id = ROMSlave_1_io_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type = ROMSlave_1_io_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type = ROMSlave_1_io_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data = ROMSlave_1_io_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready = BRAMSlave_1_io_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_valid = BRAMSlave_1_io_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat = BRAMSlave_1_io_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id = BRAMSlave_1_io_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id = BRAMSlave_1_io_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type = BRAMSlave_1_io_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type = BRAMSlave_1_io_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data = BRAMSlave_1_io_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready = PLIC_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_valid = PLIC_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat = PLIC_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id = PLIC_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id = PLIC_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type = PLIC_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type = PLIC_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data = PLIC_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_4_acquire_ready = PRCI_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_valid = PRCI_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_addr_beat = PRCI_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_client_xact_id = PRCI_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_manager_xact_id = PRCI_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_is_builtin_type = PRCI_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_g_type = PRCI_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_data = PRCI_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_5_acquire_ready = NastiIOTileLinkIOConverter_1_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_5_grant_valid = NastiIOTileLinkIOConverter_1_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_addr_beat = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_client_xact_id = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_manager_xact_id = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_is_builtin_type = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_g_type = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_5_grant_bits_data = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_data;
  assign PLIC_1_clk = clk;
  assign PLIC_1_reset = reset;
  assign PLIC_1_io_devices_0_valid = LevelGateway_2_io_plic_valid;
  assign PLIC_1_io_devices_1_valid = LevelGateway_1_1_io_plic_valid;
  assign PLIC_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid;
  assign PLIC_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block;
  assign PLIC_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id;
  assign PLIC_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat;
  assign PLIC_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type;
  assign PLIC_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type;
  assign PLIC_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union;
  assign PLIC_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data;
  assign PLIC_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_3_grant_ready;
  assign LevelGateway_2_clk = clk;
  assign LevelGateway_2_reset = reset;
  assign LevelGateway_2_io_interrupt = io_interrupts_0;
  assign LevelGateway_2_io_plic_ready = PLIC_1_io_devices_0_ready;
  assign LevelGateway_2_io_plic_complete = PLIC_1_io_devices_0_complete;
  assign LevelGateway_1_1_clk = clk;
  assign LevelGateway_1_1_reset = reset;
  assign LevelGateway_1_1_io_interrupt = io_interrupts_1;
  assign LevelGateway_1_1_io_plic_ready = PLIC_1_io_devices_1_ready;
  assign LevelGateway_1_1_io_plic_complete = PLIC_1_io_devices_1_complete;
  assign DebugModule_1_clk = clk;
  assign DebugModule_1_reset = reset;
  assign DebugModule_1_io_db_req_valid = io_debugBus_req_valid;
  assign DebugModule_1_io_db_req_bits_addr = io_debugBus_req_bits_addr;
  assign DebugModule_1_io_db_req_bits_op = io_debugBus_req_bits_op;
  assign DebugModule_1_io_db_req_bits_data = io_debugBus_req_bits_data;
  assign DebugModule_1_io_db_resp_ready = io_debugBus_resp_ready;
  assign DebugModule_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid;
  assign DebugModule_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block;
  assign DebugModule_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id;
  assign DebugModule_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat;
  assign DebugModule_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type;
  assign DebugModule_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type;
  assign DebugModule_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union;
  assign DebugModule_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data;
  assign DebugModule_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_0_grant_ready;
  assign PRCI_1_clk = clk;
  assign PRCI_1_reset = reset;
  assign PRCI_1_io_interrupts_0_meip = PLIC_1_io_harts_0;
  assign PRCI_1_io_interrupts_0_seip = PLIC_1_io_harts_1;
  assign PRCI_1_io_interrupts_0_debug = DebugModule_1_io_debugInterrupts_0;
  assign PRCI_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_4_acquire_valid;
  assign PRCI_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_block;
  assign PRCI_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_client_xact_id;
  assign PRCI_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_beat;
  assign PRCI_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_is_builtin_type;
  assign PRCI_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_a_type;
  assign PRCI_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_union;
  assign PRCI_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_data;
  assign PRCI_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_4_grant_ready;
  assign PRCI_1_io_rtcTick = T_8788;
  assign T_8788 = T_8786 == 7'h63;
  assign GEN_1 = {{6'd0}, 1'h1};
  assign T_8790 = T_8786 + GEN_1;
  assign T_8791 = T_8790[6:0];
  assign GEN_0 = T_8788 ? {{6'd0}, 1'h0} : T_8791;
  assign ROMSlave_1_clk = clk;
  assign ROMSlave_1_reset = reset;
  assign ROMSlave_1_io_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid;
  assign ROMSlave_1_io_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block;
  assign ROMSlave_1_io_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id;
  assign ROMSlave_1_io_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat;
  assign ROMSlave_1_io_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type;
  assign ROMSlave_1_io_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type;
  assign ROMSlave_1_io_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union;
  assign ROMSlave_1_io_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data;
  assign ROMSlave_1_io_grant_ready = TileLinkRecursiveInterconnect_2_io_out_1_grant_ready;
  assign BRAMSlave_1_clk = clk;
  assign BRAMSlave_1_reset = reset;
  assign BRAMSlave_1_io_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid;
  assign BRAMSlave_1_io_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block;
  assign BRAMSlave_1_io_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id;
  assign BRAMSlave_1_io_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat;
  assign BRAMSlave_1_io_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type;
  assign BRAMSlave_1_io_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type;
  assign BRAMSlave_1_io_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union;
  assign BRAMSlave_1_io_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data;
  assign BRAMSlave_1_io_grant_ready = TileLinkRecursiveInterconnect_2_io_out_2_grant_ready;
  assign NastiIOTileLinkIOConverter_1_1_clk = clk;
  assign NastiIOTileLinkIOConverter_1_1_reset = reset;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_5_acquire_valid;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_addr_block;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_client_xact_id;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_addr_beat;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_is_builtin_type;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_a_type;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_union;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_5_acquire_bits_data;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_5_grant_ready;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_aw_ready = Queue_24_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_w_ready = Queue_25_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_b_valid = Queue_27_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_resp = Queue_27_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_id = Queue_27_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_user = Queue_27_1_io_deq_bits_user;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_ar_ready = Queue_23_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_valid = Queue_26_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_resp = Queue_26_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_data = Queue_26_1_io_deq_bits_data;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_last = Queue_26_1_io_deq_bits_last;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_id = Queue_26_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_user = Queue_26_1_io_deq_bits_user;
  assign Queue_23_1_clk = clk;
  assign Queue_23_1_reset = reset;
  assign Queue_23_1_io_enq_valid = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_valid;
  assign Queue_23_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_addr;
  assign Queue_23_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_len;
  assign Queue_23_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_size;
  assign Queue_23_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_burst;
  assign Queue_23_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_lock;
  assign Queue_23_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_cache;
  assign Queue_23_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_prot;
  assign Queue_23_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_qos;
  assign Queue_23_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_region;
  assign Queue_23_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_id;
  assign Queue_23_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_user;
  assign Queue_23_1_io_deq_ready = io_mmio_axi_0_ar_ready;
  assign Queue_24_1_clk = clk;
  assign Queue_24_1_reset = reset;
  assign Queue_24_1_io_enq_valid = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_valid;
  assign Queue_24_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_addr;
  assign Queue_24_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_len;
  assign Queue_24_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_size;
  assign Queue_24_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_burst;
  assign Queue_24_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_lock;
  assign Queue_24_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_cache;
  assign Queue_24_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_prot;
  assign Queue_24_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_qos;
  assign Queue_24_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_region;
  assign Queue_24_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_id;
  assign Queue_24_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_user;
  assign Queue_24_1_io_deq_ready = io_mmio_axi_0_aw_ready;
  assign Queue_25_1_clk = clk;
  assign Queue_25_1_reset = reset;
  assign Queue_25_1_io_enq_valid = NastiIOTileLinkIOConverter_1_1_io_nasti_w_valid;
  assign Queue_25_1_io_enq_bits_data = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_data;
  assign Queue_25_1_io_enq_bits_last = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_last;
  assign Queue_25_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_id;
  assign Queue_25_1_io_enq_bits_strb = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_strb;
  assign Queue_25_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_user;
  assign Queue_25_1_io_deq_ready = io_mmio_axi_0_w_ready;
  assign Queue_26_1_clk = clk;
  assign Queue_26_1_reset = reset;
  assign Queue_26_1_io_enq_valid = io_mmio_axi_0_r_valid;
  assign Queue_26_1_io_enq_bits_resp = io_mmio_axi_0_r_bits_resp;
  assign Queue_26_1_io_enq_bits_data = io_mmio_axi_0_r_bits_data;
  assign Queue_26_1_io_enq_bits_last = io_mmio_axi_0_r_bits_last;
  assign Queue_26_1_io_enq_bits_id = io_mmio_axi_0_r_bits_id;
  assign Queue_26_1_io_enq_bits_user = io_mmio_axi_0_r_bits_user;
  assign Queue_26_1_io_deq_ready = NastiIOTileLinkIOConverter_1_1_io_nasti_r_ready;
  assign Queue_27_1_clk = clk;
  assign Queue_27_1_reset = reset;
  assign Queue_27_1_io_enq_valid = io_mmio_axi_0_b_valid;
  assign Queue_27_1_io_enq_bits_resp = io_mmio_axi_0_b_bits_resp;
  assign Queue_27_1_io_enq_bits_id = io_mmio_axi_0_b_bits_id;
  assign Queue_27_1_io_enq_bits_user = io_mmio_axi_0_b_bits_user;
  assign Queue_27_1_io_deq_ready = NastiIOTileLinkIOConverter_1_1_io_nasti_b_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_2 = {1{$random}};
  T_8786 = GEN_2[6:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_8786 <= 7'h0;
    end else begin
      if(T_8788) begin
        T_8786 <= {{6'd0}, 1'h0};
      end else begin
        T_8786 <= T_8791;
      end
    end
  end
endmodule
module Top(
  input   clk,
  input   reset,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  input   io_interrupts_0,
  input   io_interrupts_1,
  input   io_mmio_axi_0_aw_ready,
  output  io_mmio_axi_0_aw_valid,
  output [31:0] io_mmio_axi_0_aw_bits_addr,
  output [7:0] io_mmio_axi_0_aw_bits_len,
  output [2:0] io_mmio_axi_0_aw_bits_size,
  output [1:0] io_mmio_axi_0_aw_bits_burst,
  output  io_mmio_axi_0_aw_bits_lock,
  output [3:0] io_mmio_axi_0_aw_bits_cache,
  output [2:0] io_mmio_axi_0_aw_bits_prot,
  output [3:0] io_mmio_axi_0_aw_bits_qos,
  output [3:0] io_mmio_axi_0_aw_bits_region,
  output [4:0] io_mmio_axi_0_aw_bits_id,
  output  io_mmio_axi_0_aw_bits_user,
  input   io_mmio_axi_0_w_ready,
  output  io_mmio_axi_0_w_valid,
  output [63:0] io_mmio_axi_0_w_bits_data,
  output  io_mmio_axi_0_w_bits_last,
  output [4:0] io_mmio_axi_0_w_bits_id,
  output [7:0] io_mmio_axi_0_w_bits_strb,
  output  io_mmio_axi_0_w_bits_user,
  output  io_mmio_axi_0_b_ready,
  input   io_mmio_axi_0_b_valid,
  input  [1:0] io_mmio_axi_0_b_bits_resp,
  input  [4:0] io_mmio_axi_0_b_bits_id,
  input   io_mmio_axi_0_b_bits_user,
  input   io_mmio_axi_0_ar_ready,
  output  io_mmio_axi_0_ar_valid,
  output [31:0] io_mmio_axi_0_ar_bits_addr,
  output [7:0] io_mmio_axi_0_ar_bits_len,
  output [2:0] io_mmio_axi_0_ar_bits_size,
  output [1:0] io_mmio_axi_0_ar_bits_burst,
  output  io_mmio_axi_0_ar_bits_lock,
  output [3:0] io_mmio_axi_0_ar_bits_cache,
  output [2:0] io_mmio_axi_0_ar_bits_prot,
  output [3:0] io_mmio_axi_0_ar_bits_qos,
  output [3:0] io_mmio_axi_0_ar_bits_region,
  output [4:0] io_mmio_axi_0_ar_bits_id,
  output  io_mmio_axi_0_ar_bits_user,
  output  io_mmio_axi_0_r_ready,
  input   io_mmio_axi_0_r_valid,
  input  [1:0] io_mmio_axi_0_r_bits_resp,
  input  [63:0] io_mmio_axi_0_r_bits_data,
  input   io_mmio_axi_0_r_bits_last,
  input  [4:0] io_mmio_axi_0_r_bits_id,
  input   io_mmio_axi_0_r_bits_user,
  output  io_debug_req_ready,
  input   io_debug_req_valid,
  input  [4:0] io_debug_req_bits_addr,
  input  [1:0] io_debug_req_bits_op,
  input  [33:0] io_debug_req_bits_data,
  input   io_debug_resp_ready,
  output  io_debug_resp_valid,
  output [1:0] io_debug_resp_bits_resp,
  output [33:0] io_debug_resp_bits_data
);
  wire  tileResets_0;
  wire  RocketTile_1_clk;
  wire  RocketTile_1_reset;
  wire  RocketTile_1_io_cached_0_acquire_ready;
  wire  RocketTile_1_io_cached_0_acquire_valid;
  wire [25:0] RocketTile_1_io_cached_0_acquire_bits_addr_block;
  wire [1:0] RocketTile_1_io_cached_0_acquire_bits_client_xact_id;
  wire [2:0] RocketTile_1_io_cached_0_acquire_bits_addr_beat;
  wire  RocketTile_1_io_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] RocketTile_1_io_cached_0_acquire_bits_a_type;
  wire [11:0] RocketTile_1_io_cached_0_acquire_bits_union;
  wire [63:0] RocketTile_1_io_cached_0_acquire_bits_data;
  wire  RocketTile_1_io_cached_0_probe_ready;
  wire  RocketTile_1_io_cached_0_probe_valid;
  wire [25:0] RocketTile_1_io_cached_0_probe_bits_addr_block;
  wire [1:0] RocketTile_1_io_cached_0_probe_bits_p_type;
  wire  RocketTile_1_io_cached_0_release_ready;
  wire  RocketTile_1_io_cached_0_release_valid;
  wire [2:0] RocketTile_1_io_cached_0_release_bits_addr_beat;
  wire [25:0] RocketTile_1_io_cached_0_release_bits_addr_block;
  wire [1:0] RocketTile_1_io_cached_0_release_bits_client_xact_id;
  wire  RocketTile_1_io_cached_0_release_bits_voluntary;
  wire [2:0] RocketTile_1_io_cached_0_release_bits_r_type;
  wire [63:0] RocketTile_1_io_cached_0_release_bits_data;
  wire  RocketTile_1_io_cached_0_grant_ready;
  wire  RocketTile_1_io_cached_0_grant_valid;
  wire [2:0] RocketTile_1_io_cached_0_grant_bits_addr_beat;
  wire [1:0] RocketTile_1_io_cached_0_grant_bits_client_xact_id;
  wire [2:0] RocketTile_1_io_cached_0_grant_bits_manager_xact_id;
  wire  RocketTile_1_io_cached_0_grant_bits_is_builtin_type;
  wire [3:0] RocketTile_1_io_cached_0_grant_bits_g_type;
  wire [63:0] RocketTile_1_io_cached_0_grant_bits_data;
  wire  RocketTile_1_io_cached_0_grant_bits_manager_id;
  wire  RocketTile_1_io_cached_0_finish_ready;
  wire  RocketTile_1_io_cached_0_finish_valid;
  wire [2:0] RocketTile_1_io_cached_0_finish_bits_manager_xact_id;
  wire  RocketTile_1_io_cached_0_finish_bits_manager_id;
  wire  RocketTile_1_io_uncached_0_acquire_ready;
  wire  RocketTile_1_io_uncached_0_acquire_valid;
  wire [25:0] RocketTile_1_io_uncached_0_acquire_bits_addr_block;
  wire [1:0] RocketTile_1_io_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] RocketTile_1_io_uncached_0_acquire_bits_addr_beat;
  wire  RocketTile_1_io_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] RocketTile_1_io_uncached_0_acquire_bits_a_type;
  wire [11:0] RocketTile_1_io_uncached_0_acquire_bits_union;
  wire [63:0] RocketTile_1_io_uncached_0_acquire_bits_data;
  wire  RocketTile_1_io_uncached_0_grant_ready;
  wire  RocketTile_1_io_uncached_0_grant_valid;
  wire [2:0] RocketTile_1_io_uncached_0_grant_bits_addr_beat;
  wire [1:0] RocketTile_1_io_uncached_0_grant_bits_client_xact_id;
  wire [2:0] RocketTile_1_io_uncached_0_grant_bits_manager_xact_id;
  wire  RocketTile_1_io_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] RocketTile_1_io_uncached_0_grant_bits_g_type;
  wire [63:0] RocketTile_1_io_uncached_0_grant_bits_data;
  wire  RocketTile_1_io_prci_reset;
  wire  RocketTile_1_io_prci_id;
  wire  RocketTile_1_io_prci_interrupts_meip;
  wire  RocketTile_1_io_prci_interrupts_seip;
  wire  RocketTile_1_io_prci_interrupts_debug;
  wire  RocketTile_1_io_prci_interrupts_mtip;
  wire  RocketTile_1_io_prci_interrupts_msip;
  wire  uncore_clk;
  wire  uncore_reset;
  wire  uncore_io_mem_axi_0_aw_ready;
  wire  uncore_io_mem_axi_0_aw_valid;
  wire [31:0] uncore_io_mem_axi_0_aw_bits_addr;
  wire [7:0] uncore_io_mem_axi_0_aw_bits_len;
  wire [2:0] uncore_io_mem_axi_0_aw_bits_size;
  wire [1:0] uncore_io_mem_axi_0_aw_bits_burst;
  wire  uncore_io_mem_axi_0_aw_bits_lock;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_cache;
  wire [2:0] uncore_io_mem_axi_0_aw_bits_prot;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_qos;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_region;
  wire [4:0] uncore_io_mem_axi_0_aw_bits_id;
  wire  uncore_io_mem_axi_0_aw_bits_user;
  wire  uncore_io_mem_axi_0_w_ready;
  wire  uncore_io_mem_axi_0_w_valid;
  wire [63:0] uncore_io_mem_axi_0_w_bits_data;
  wire  uncore_io_mem_axi_0_w_bits_last;
  wire [4:0] uncore_io_mem_axi_0_w_bits_id;
  wire [7:0] uncore_io_mem_axi_0_w_bits_strb;
  wire  uncore_io_mem_axi_0_w_bits_user;
  wire  uncore_io_mem_axi_0_b_ready;
  wire  uncore_io_mem_axi_0_b_valid;
  wire [1:0] uncore_io_mem_axi_0_b_bits_resp;
  wire [4:0] uncore_io_mem_axi_0_b_bits_id;
  wire  uncore_io_mem_axi_0_b_bits_user;
  wire  uncore_io_mem_axi_0_ar_ready;
  wire  uncore_io_mem_axi_0_ar_valid;
  wire [31:0] uncore_io_mem_axi_0_ar_bits_addr;
  wire [7:0] uncore_io_mem_axi_0_ar_bits_len;
  wire [2:0] uncore_io_mem_axi_0_ar_bits_size;
  wire [1:0] uncore_io_mem_axi_0_ar_bits_burst;
  wire  uncore_io_mem_axi_0_ar_bits_lock;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_cache;
  wire [2:0] uncore_io_mem_axi_0_ar_bits_prot;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_qos;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_region;
  wire [4:0] uncore_io_mem_axi_0_ar_bits_id;
  wire  uncore_io_mem_axi_0_ar_bits_user;
  wire  uncore_io_mem_axi_0_r_ready;
  wire  uncore_io_mem_axi_0_r_valid;
  wire [1:0] uncore_io_mem_axi_0_r_bits_resp;
  wire [63:0] uncore_io_mem_axi_0_r_bits_data;
  wire  uncore_io_mem_axi_0_r_bits_last;
  wire [4:0] uncore_io_mem_axi_0_r_bits_id;
  wire  uncore_io_mem_axi_0_r_bits_user;
  wire  uncore_io_tiles_cached_0_acquire_ready;
  wire  uncore_io_tiles_cached_0_acquire_valid;
  wire [25:0] uncore_io_tiles_cached_0_acquire_bits_addr_block;
  wire [1:0] uncore_io_tiles_cached_0_acquire_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_cached_0_acquire_bits_addr_beat;
  wire  uncore_io_tiles_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] uncore_io_tiles_cached_0_acquire_bits_a_type;
  wire [11:0] uncore_io_tiles_cached_0_acquire_bits_union;
  wire [63:0] uncore_io_tiles_cached_0_acquire_bits_data;
  wire  uncore_io_tiles_cached_0_probe_ready;
  wire  uncore_io_tiles_cached_0_probe_valid;
  wire [25:0] uncore_io_tiles_cached_0_probe_bits_addr_block;
  wire [1:0] uncore_io_tiles_cached_0_probe_bits_p_type;
  wire  uncore_io_tiles_cached_0_release_ready;
  wire  uncore_io_tiles_cached_0_release_valid;
  wire [2:0] uncore_io_tiles_cached_0_release_bits_addr_beat;
  wire [25:0] uncore_io_tiles_cached_0_release_bits_addr_block;
  wire [1:0] uncore_io_tiles_cached_0_release_bits_client_xact_id;
  wire  uncore_io_tiles_cached_0_release_bits_voluntary;
  wire [2:0] uncore_io_tiles_cached_0_release_bits_r_type;
  wire [63:0] uncore_io_tiles_cached_0_release_bits_data;
  wire  uncore_io_tiles_cached_0_grant_ready;
  wire  uncore_io_tiles_cached_0_grant_valid;
  wire [2:0] uncore_io_tiles_cached_0_grant_bits_addr_beat;
  wire [1:0] uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire  uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire [3:0] uncore_io_tiles_cached_0_grant_bits_g_type;
  wire [63:0] uncore_io_tiles_cached_0_grant_bits_data;
  wire  uncore_io_tiles_cached_0_grant_bits_manager_id;
  wire  uncore_io_tiles_cached_0_finish_ready;
  wire  uncore_io_tiles_cached_0_finish_valid;
  wire [2:0] uncore_io_tiles_cached_0_finish_bits_manager_xact_id;
  wire  uncore_io_tiles_cached_0_finish_bits_manager_id;
  wire  uncore_io_tiles_uncached_0_acquire_ready;
  wire  uncore_io_tiles_uncached_0_acquire_valid;
  wire [25:0] uncore_io_tiles_uncached_0_acquire_bits_addr_block;
  wire [1:0] uncore_io_tiles_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_uncached_0_acquire_bits_addr_beat;
  wire  uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] uncore_io_tiles_uncached_0_acquire_bits_a_type;
  wire [11:0] uncore_io_tiles_uncached_0_acquire_bits_union;
  wire [63:0] uncore_io_tiles_uncached_0_acquire_bits_data;
  wire  uncore_io_tiles_uncached_0_grant_ready;
  wire  uncore_io_tiles_uncached_0_grant_valid;
  wire [2:0] uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  wire [1:0] uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire  uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] uncore_io_tiles_uncached_0_grant_bits_g_type;
  wire [63:0] uncore_io_tiles_uncached_0_grant_bits_data;
  wire  uncore_io_prci_0_reset;
  wire  uncore_io_prci_0_id;
  wire  uncore_io_prci_0_interrupts_meip;
  wire  uncore_io_prci_0_interrupts_seip;
  wire  uncore_io_prci_0_interrupts_debug;
  wire  uncore_io_prci_0_interrupts_mtip;
  wire  uncore_io_prci_0_interrupts_msip;
  wire  uncore_io_mmio_axi_0_aw_ready;
  wire  uncore_io_mmio_axi_0_aw_valid;
  wire [31:0] uncore_io_mmio_axi_0_aw_bits_addr;
  wire [7:0] uncore_io_mmio_axi_0_aw_bits_len;
  wire [2:0] uncore_io_mmio_axi_0_aw_bits_size;
  wire [1:0] uncore_io_mmio_axi_0_aw_bits_burst;
  wire  uncore_io_mmio_axi_0_aw_bits_lock;
  wire [3:0] uncore_io_mmio_axi_0_aw_bits_cache;
  wire [2:0] uncore_io_mmio_axi_0_aw_bits_prot;
  wire [3:0] uncore_io_mmio_axi_0_aw_bits_qos;
  wire [3:0] uncore_io_mmio_axi_0_aw_bits_region;
  wire [4:0] uncore_io_mmio_axi_0_aw_bits_id;
  wire  uncore_io_mmio_axi_0_aw_bits_user;
  wire  uncore_io_mmio_axi_0_w_ready;
  wire  uncore_io_mmio_axi_0_w_valid;
  wire [63:0] uncore_io_mmio_axi_0_w_bits_data;
  wire  uncore_io_mmio_axi_0_w_bits_last;
  wire [4:0] uncore_io_mmio_axi_0_w_bits_id;
  wire [7:0] uncore_io_mmio_axi_0_w_bits_strb;
  wire  uncore_io_mmio_axi_0_w_bits_user;
  wire  uncore_io_mmio_axi_0_b_ready;
  wire  uncore_io_mmio_axi_0_b_valid;
  wire [1:0] uncore_io_mmio_axi_0_b_bits_resp;
  wire [4:0] uncore_io_mmio_axi_0_b_bits_id;
  wire  uncore_io_mmio_axi_0_b_bits_user;
  wire  uncore_io_mmio_axi_0_ar_ready;
  wire  uncore_io_mmio_axi_0_ar_valid;
  wire [31:0] uncore_io_mmio_axi_0_ar_bits_addr;
  wire [7:0] uncore_io_mmio_axi_0_ar_bits_len;
  wire [2:0] uncore_io_mmio_axi_0_ar_bits_size;
  wire [1:0] uncore_io_mmio_axi_0_ar_bits_burst;
  wire  uncore_io_mmio_axi_0_ar_bits_lock;
  wire [3:0] uncore_io_mmio_axi_0_ar_bits_cache;
  wire [2:0] uncore_io_mmio_axi_0_ar_bits_prot;
  wire [3:0] uncore_io_mmio_axi_0_ar_bits_qos;
  wire [3:0] uncore_io_mmio_axi_0_ar_bits_region;
  wire [4:0] uncore_io_mmio_axi_0_ar_bits_id;
  wire  uncore_io_mmio_axi_0_ar_bits_user;
  wire  uncore_io_mmio_axi_0_r_ready;
  wire  uncore_io_mmio_axi_0_r_valid;
  wire [1:0] uncore_io_mmio_axi_0_r_bits_resp;
  wire [63:0] uncore_io_mmio_axi_0_r_bits_data;
  wire  uncore_io_mmio_axi_0_r_bits_last;
  wire [4:0] uncore_io_mmio_axi_0_r_bits_id;
  wire  uncore_io_mmio_axi_0_r_bits_user;
  wire  uncore_io_interrupts_0;
  wire  uncore_io_interrupts_1;
  wire  uncore_io_debugBus_req_ready;
  wire  uncore_io_debugBus_req_valid;
  wire [4:0] uncore_io_debugBus_req_bits_addr;
  wire [1:0] uncore_io_debugBus_req_bits_op;
  wire [33:0] uncore_io_debugBus_req_bits_data;
  wire  uncore_io_debugBus_resp_ready;
  wire  uncore_io_debugBus_resp_valid;
  wire [1:0] uncore_io_debugBus_resp_bits_resp;
  wire [33:0] uncore_io_debugBus_resp_bits_data;
  RocketTile RocketTile_1 (
    .clk(RocketTile_1_clk),
    .reset(RocketTile_1_reset),
    .io_cached_0_acquire_ready(RocketTile_1_io_cached_0_acquire_ready),
    .io_cached_0_acquire_valid(RocketTile_1_io_cached_0_acquire_valid),
    .io_cached_0_acquire_bits_addr_block(RocketTile_1_io_cached_0_acquire_bits_addr_block),
    .io_cached_0_acquire_bits_client_xact_id(RocketTile_1_io_cached_0_acquire_bits_client_xact_id),
    .io_cached_0_acquire_bits_addr_beat(RocketTile_1_io_cached_0_acquire_bits_addr_beat),
    .io_cached_0_acquire_bits_is_builtin_type(RocketTile_1_io_cached_0_acquire_bits_is_builtin_type),
    .io_cached_0_acquire_bits_a_type(RocketTile_1_io_cached_0_acquire_bits_a_type),
    .io_cached_0_acquire_bits_union(RocketTile_1_io_cached_0_acquire_bits_union),
    .io_cached_0_acquire_bits_data(RocketTile_1_io_cached_0_acquire_bits_data),
    .io_cached_0_probe_ready(RocketTile_1_io_cached_0_probe_ready),
    .io_cached_0_probe_valid(RocketTile_1_io_cached_0_probe_valid),
    .io_cached_0_probe_bits_addr_block(RocketTile_1_io_cached_0_probe_bits_addr_block),
    .io_cached_0_probe_bits_p_type(RocketTile_1_io_cached_0_probe_bits_p_type),
    .io_cached_0_release_ready(RocketTile_1_io_cached_0_release_ready),
    .io_cached_0_release_valid(RocketTile_1_io_cached_0_release_valid),
    .io_cached_0_release_bits_addr_beat(RocketTile_1_io_cached_0_release_bits_addr_beat),
    .io_cached_0_release_bits_addr_block(RocketTile_1_io_cached_0_release_bits_addr_block),
    .io_cached_0_release_bits_client_xact_id(RocketTile_1_io_cached_0_release_bits_client_xact_id),
    .io_cached_0_release_bits_voluntary(RocketTile_1_io_cached_0_release_bits_voluntary),
    .io_cached_0_release_bits_r_type(RocketTile_1_io_cached_0_release_bits_r_type),
    .io_cached_0_release_bits_data(RocketTile_1_io_cached_0_release_bits_data),
    .io_cached_0_grant_ready(RocketTile_1_io_cached_0_grant_ready),
    .io_cached_0_grant_valid(RocketTile_1_io_cached_0_grant_valid),
    .io_cached_0_grant_bits_addr_beat(RocketTile_1_io_cached_0_grant_bits_addr_beat),
    .io_cached_0_grant_bits_client_xact_id(RocketTile_1_io_cached_0_grant_bits_client_xact_id),
    .io_cached_0_grant_bits_manager_xact_id(RocketTile_1_io_cached_0_grant_bits_manager_xact_id),
    .io_cached_0_grant_bits_is_builtin_type(RocketTile_1_io_cached_0_grant_bits_is_builtin_type),
    .io_cached_0_grant_bits_g_type(RocketTile_1_io_cached_0_grant_bits_g_type),
    .io_cached_0_grant_bits_data(RocketTile_1_io_cached_0_grant_bits_data),
    .io_cached_0_grant_bits_manager_id(RocketTile_1_io_cached_0_grant_bits_manager_id),
    .io_cached_0_finish_ready(RocketTile_1_io_cached_0_finish_ready),
    .io_cached_0_finish_valid(RocketTile_1_io_cached_0_finish_valid),
    .io_cached_0_finish_bits_manager_xact_id(RocketTile_1_io_cached_0_finish_bits_manager_xact_id),
    .io_cached_0_finish_bits_manager_id(RocketTile_1_io_cached_0_finish_bits_manager_id),
    .io_uncached_0_acquire_ready(RocketTile_1_io_uncached_0_acquire_ready),
    .io_uncached_0_acquire_valid(RocketTile_1_io_uncached_0_acquire_valid),
    .io_uncached_0_acquire_bits_addr_block(RocketTile_1_io_uncached_0_acquire_bits_addr_block),
    .io_uncached_0_acquire_bits_client_xact_id(RocketTile_1_io_uncached_0_acquire_bits_client_xact_id),
    .io_uncached_0_acquire_bits_addr_beat(RocketTile_1_io_uncached_0_acquire_bits_addr_beat),
    .io_uncached_0_acquire_bits_is_builtin_type(RocketTile_1_io_uncached_0_acquire_bits_is_builtin_type),
    .io_uncached_0_acquire_bits_a_type(RocketTile_1_io_uncached_0_acquire_bits_a_type),
    .io_uncached_0_acquire_bits_union(RocketTile_1_io_uncached_0_acquire_bits_union),
    .io_uncached_0_acquire_bits_data(RocketTile_1_io_uncached_0_acquire_bits_data),
    .io_uncached_0_grant_ready(RocketTile_1_io_uncached_0_grant_ready),
    .io_uncached_0_grant_valid(RocketTile_1_io_uncached_0_grant_valid),
    .io_uncached_0_grant_bits_addr_beat(RocketTile_1_io_uncached_0_grant_bits_addr_beat),
    .io_uncached_0_grant_bits_client_xact_id(RocketTile_1_io_uncached_0_grant_bits_client_xact_id),
    .io_uncached_0_grant_bits_manager_xact_id(RocketTile_1_io_uncached_0_grant_bits_manager_xact_id),
    .io_uncached_0_grant_bits_is_builtin_type(RocketTile_1_io_uncached_0_grant_bits_is_builtin_type),
    .io_uncached_0_grant_bits_g_type(RocketTile_1_io_uncached_0_grant_bits_g_type),
    .io_uncached_0_grant_bits_data(RocketTile_1_io_uncached_0_grant_bits_data),
    .io_prci_reset(RocketTile_1_io_prci_reset),
    .io_prci_id(RocketTile_1_io_prci_id),
    .io_prci_interrupts_meip(RocketTile_1_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(RocketTile_1_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(RocketTile_1_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(RocketTile_1_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(RocketTile_1_io_prci_interrupts_msip)
  );
  Uncore uncore (
    .clk(uncore_clk),
    .reset(uncore_reset),
    .io_mem_axi_0_aw_ready(uncore_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(uncore_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(uncore_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(uncore_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(uncore_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(uncore_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(uncore_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(uncore_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(uncore_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(uncore_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(uncore_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(uncore_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(uncore_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(uncore_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(uncore_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(uncore_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(uncore_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(uncore_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(uncore_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(uncore_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(uncore_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(uncore_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(uncore_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(uncore_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(uncore_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(uncore_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(uncore_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(uncore_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(uncore_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(uncore_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(uncore_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(uncore_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(uncore_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(uncore_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(uncore_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(uncore_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(uncore_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(uncore_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(uncore_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(uncore_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(uncore_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(uncore_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(uncore_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(uncore_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(uncore_io_mem_axi_0_r_bits_user),
    .io_tiles_cached_0_acquire_ready(uncore_io_tiles_cached_0_acquire_ready),
    .io_tiles_cached_0_acquire_valid(uncore_io_tiles_cached_0_acquire_valid),
    .io_tiles_cached_0_acquire_bits_addr_block(uncore_io_tiles_cached_0_acquire_bits_addr_block),
    .io_tiles_cached_0_acquire_bits_client_xact_id(uncore_io_tiles_cached_0_acquire_bits_client_xact_id),
    .io_tiles_cached_0_acquire_bits_addr_beat(uncore_io_tiles_cached_0_acquire_bits_addr_beat),
    .io_tiles_cached_0_acquire_bits_is_builtin_type(uncore_io_tiles_cached_0_acquire_bits_is_builtin_type),
    .io_tiles_cached_0_acquire_bits_a_type(uncore_io_tiles_cached_0_acquire_bits_a_type),
    .io_tiles_cached_0_acquire_bits_union(uncore_io_tiles_cached_0_acquire_bits_union),
    .io_tiles_cached_0_acquire_bits_data(uncore_io_tiles_cached_0_acquire_bits_data),
    .io_tiles_cached_0_probe_ready(uncore_io_tiles_cached_0_probe_ready),
    .io_tiles_cached_0_probe_valid(uncore_io_tiles_cached_0_probe_valid),
    .io_tiles_cached_0_probe_bits_addr_block(uncore_io_tiles_cached_0_probe_bits_addr_block),
    .io_tiles_cached_0_probe_bits_p_type(uncore_io_tiles_cached_0_probe_bits_p_type),
    .io_tiles_cached_0_release_ready(uncore_io_tiles_cached_0_release_ready),
    .io_tiles_cached_0_release_valid(uncore_io_tiles_cached_0_release_valid),
    .io_tiles_cached_0_release_bits_addr_beat(uncore_io_tiles_cached_0_release_bits_addr_beat),
    .io_tiles_cached_0_release_bits_addr_block(uncore_io_tiles_cached_0_release_bits_addr_block),
    .io_tiles_cached_0_release_bits_client_xact_id(uncore_io_tiles_cached_0_release_bits_client_xact_id),
    .io_tiles_cached_0_release_bits_voluntary(uncore_io_tiles_cached_0_release_bits_voluntary),
    .io_tiles_cached_0_release_bits_r_type(uncore_io_tiles_cached_0_release_bits_r_type),
    .io_tiles_cached_0_release_bits_data(uncore_io_tiles_cached_0_release_bits_data),
    .io_tiles_cached_0_grant_ready(uncore_io_tiles_cached_0_grant_ready),
    .io_tiles_cached_0_grant_valid(uncore_io_tiles_cached_0_grant_valid),
    .io_tiles_cached_0_grant_bits_addr_beat(uncore_io_tiles_cached_0_grant_bits_addr_beat),
    .io_tiles_cached_0_grant_bits_client_xact_id(uncore_io_tiles_cached_0_grant_bits_client_xact_id),
    .io_tiles_cached_0_grant_bits_manager_xact_id(uncore_io_tiles_cached_0_grant_bits_manager_xact_id),
    .io_tiles_cached_0_grant_bits_is_builtin_type(uncore_io_tiles_cached_0_grant_bits_is_builtin_type),
    .io_tiles_cached_0_grant_bits_g_type(uncore_io_tiles_cached_0_grant_bits_g_type),
    .io_tiles_cached_0_grant_bits_data(uncore_io_tiles_cached_0_grant_bits_data),
    .io_tiles_cached_0_grant_bits_manager_id(uncore_io_tiles_cached_0_grant_bits_manager_id),
    .io_tiles_cached_0_finish_ready(uncore_io_tiles_cached_0_finish_ready),
    .io_tiles_cached_0_finish_valid(uncore_io_tiles_cached_0_finish_valid),
    .io_tiles_cached_0_finish_bits_manager_xact_id(uncore_io_tiles_cached_0_finish_bits_manager_xact_id),
    .io_tiles_cached_0_finish_bits_manager_id(uncore_io_tiles_cached_0_finish_bits_manager_id),
    .io_tiles_uncached_0_acquire_ready(uncore_io_tiles_uncached_0_acquire_ready),
    .io_tiles_uncached_0_acquire_valid(uncore_io_tiles_uncached_0_acquire_valid),
    .io_tiles_uncached_0_acquire_bits_addr_block(uncore_io_tiles_uncached_0_acquire_bits_addr_block),
    .io_tiles_uncached_0_acquire_bits_client_xact_id(uncore_io_tiles_uncached_0_acquire_bits_client_xact_id),
    .io_tiles_uncached_0_acquire_bits_addr_beat(uncore_io_tiles_uncached_0_acquire_bits_addr_beat),
    .io_tiles_uncached_0_acquire_bits_is_builtin_type(uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type),
    .io_tiles_uncached_0_acquire_bits_a_type(uncore_io_tiles_uncached_0_acquire_bits_a_type),
    .io_tiles_uncached_0_acquire_bits_union(uncore_io_tiles_uncached_0_acquire_bits_union),
    .io_tiles_uncached_0_acquire_bits_data(uncore_io_tiles_uncached_0_acquire_bits_data),
    .io_tiles_uncached_0_grant_ready(uncore_io_tiles_uncached_0_grant_ready),
    .io_tiles_uncached_0_grant_valid(uncore_io_tiles_uncached_0_grant_valid),
    .io_tiles_uncached_0_grant_bits_addr_beat(uncore_io_tiles_uncached_0_grant_bits_addr_beat),
    .io_tiles_uncached_0_grant_bits_client_xact_id(uncore_io_tiles_uncached_0_grant_bits_client_xact_id),
    .io_tiles_uncached_0_grant_bits_manager_xact_id(uncore_io_tiles_uncached_0_grant_bits_manager_xact_id),
    .io_tiles_uncached_0_grant_bits_is_builtin_type(uncore_io_tiles_uncached_0_grant_bits_is_builtin_type),
    .io_tiles_uncached_0_grant_bits_g_type(uncore_io_tiles_uncached_0_grant_bits_g_type),
    .io_tiles_uncached_0_grant_bits_data(uncore_io_tiles_uncached_0_grant_bits_data),
    .io_prci_0_reset(uncore_io_prci_0_reset),
    .io_prci_0_id(uncore_io_prci_0_id),
    .io_prci_0_interrupts_meip(uncore_io_prci_0_interrupts_meip),
    .io_prci_0_interrupts_seip(uncore_io_prci_0_interrupts_seip),
    .io_prci_0_interrupts_debug(uncore_io_prci_0_interrupts_debug),
    .io_prci_0_interrupts_mtip(uncore_io_prci_0_interrupts_mtip),
    .io_prci_0_interrupts_msip(uncore_io_prci_0_interrupts_msip),
    .io_mmio_axi_0_aw_ready(uncore_io_mmio_axi_0_aw_ready),
    .io_mmio_axi_0_aw_valid(uncore_io_mmio_axi_0_aw_valid),
    .io_mmio_axi_0_aw_bits_addr(uncore_io_mmio_axi_0_aw_bits_addr),
    .io_mmio_axi_0_aw_bits_len(uncore_io_mmio_axi_0_aw_bits_len),
    .io_mmio_axi_0_aw_bits_size(uncore_io_mmio_axi_0_aw_bits_size),
    .io_mmio_axi_0_aw_bits_burst(uncore_io_mmio_axi_0_aw_bits_burst),
    .io_mmio_axi_0_aw_bits_lock(uncore_io_mmio_axi_0_aw_bits_lock),
    .io_mmio_axi_0_aw_bits_cache(uncore_io_mmio_axi_0_aw_bits_cache),
    .io_mmio_axi_0_aw_bits_prot(uncore_io_mmio_axi_0_aw_bits_prot),
    .io_mmio_axi_0_aw_bits_qos(uncore_io_mmio_axi_0_aw_bits_qos),
    .io_mmio_axi_0_aw_bits_region(uncore_io_mmio_axi_0_aw_bits_region),
    .io_mmio_axi_0_aw_bits_id(uncore_io_mmio_axi_0_aw_bits_id),
    .io_mmio_axi_0_aw_bits_user(uncore_io_mmio_axi_0_aw_bits_user),
    .io_mmio_axi_0_w_ready(uncore_io_mmio_axi_0_w_ready),
    .io_mmio_axi_0_w_valid(uncore_io_mmio_axi_0_w_valid),
    .io_mmio_axi_0_w_bits_data(uncore_io_mmio_axi_0_w_bits_data),
    .io_mmio_axi_0_w_bits_last(uncore_io_mmio_axi_0_w_bits_last),
    .io_mmio_axi_0_w_bits_id(uncore_io_mmio_axi_0_w_bits_id),
    .io_mmio_axi_0_w_bits_strb(uncore_io_mmio_axi_0_w_bits_strb),
    .io_mmio_axi_0_w_bits_user(uncore_io_mmio_axi_0_w_bits_user),
    .io_mmio_axi_0_b_ready(uncore_io_mmio_axi_0_b_ready),
    .io_mmio_axi_0_b_valid(uncore_io_mmio_axi_0_b_valid),
    .io_mmio_axi_0_b_bits_resp(uncore_io_mmio_axi_0_b_bits_resp),
    .io_mmio_axi_0_b_bits_id(uncore_io_mmio_axi_0_b_bits_id),
    .io_mmio_axi_0_b_bits_user(uncore_io_mmio_axi_0_b_bits_user),
    .io_mmio_axi_0_ar_ready(uncore_io_mmio_axi_0_ar_ready),
    .io_mmio_axi_0_ar_valid(uncore_io_mmio_axi_0_ar_valid),
    .io_mmio_axi_0_ar_bits_addr(uncore_io_mmio_axi_0_ar_bits_addr),
    .io_mmio_axi_0_ar_bits_len(uncore_io_mmio_axi_0_ar_bits_len),
    .io_mmio_axi_0_ar_bits_size(uncore_io_mmio_axi_0_ar_bits_size),
    .io_mmio_axi_0_ar_bits_burst(uncore_io_mmio_axi_0_ar_bits_burst),
    .io_mmio_axi_0_ar_bits_lock(uncore_io_mmio_axi_0_ar_bits_lock),
    .io_mmio_axi_0_ar_bits_cache(uncore_io_mmio_axi_0_ar_bits_cache),
    .io_mmio_axi_0_ar_bits_prot(uncore_io_mmio_axi_0_ar_bits_prot),
    .io_mmio_axi_0_ar_bits_qos(uncore_io_mmio_axi_0_ar_bits_qos),
    .io_mmio_axi_0_ar_bits_region(uncore_io_mmio_axi_0_ar_bits_region),
    .io_mmio_axi_0_ar_bits_id(uncore_io_mmio_axi_0_ar_bits_id),
    .io_mmio_axi_0_ar_bits_user(uncore_io_mmio_axi_0_ar_bits_user),
    .io_mmio_axi_0_r_ready(uncore_io_mmio_axi_0_r_ready),
    .io_mmio_axi_0_r_valid(uncore_io_mmio_axi_0_r_valid),
    .io_mmio_axi_0_r_bits_resp(uncore_io_mmio_axi_0_r_bits_resp),
    .io_mmio_axi_0_r_bits_data(uncore_io_mmio_axi_0_r_bits_data),
    .io_mmio_axi_0_r_bits_last(uncore_io_mmio_axi_0_r_bits_last),
    .io_mmio_axi_0_r_bits_id(uncore_io_mmio_axi_0_r_bits_id),
    .io_mmio_axi_0_r_bits_user(uncore_io_mmio_axi_0_r_bits_user),
    .io_interrupts_0(uncore_io_interrupts_0),
    .io_interrupts_1(uncore_io_interrupts_1),
    .io_debugBus_req_ready(uncore_io_debugBus_req_ready),
    .io_debugBus_req_valid(uncore_io_debugBus_req_valid),
    .io_debugBus_req_bits_addr(uncore_io_debugBus_req_bits_addr),
    .io_debugBus_req_bits_op(uncore_io_debugBus_req_bits_op),
    .io_debugBus_req_bits_data(uncore_io_debugBus_req_bits_data),
    .io_debugBus_resp_ready(uncore_io_debugBus_resp_ready),
    .io_debugBus_resp_valid(uncore_io_debugBus_resp_valid),
    .io_debugBus_resp_bits_resp(uncore_io_debugBus_resp_bits_resp),
    .io_debugBus_resp_bits_data(uncore_io_debugBus_resp_bits_data)
  );
  assign io_mem_axi_0_aw_valid = uncore_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = uncore_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = uncore_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = uncore_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = uncore_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = uncore_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = uncore_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = uncore_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = uncore_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = uncore_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = uncore_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = uncore_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = uncore_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = uncore_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = uncore_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = uncore_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = uncore_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = uncore_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = uncore_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = uncore_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = uncore_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = uncore_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = uncore_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = uncore_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = uncore_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = uncore_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = uncore_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = uncore_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = uncore_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = uncore_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = uncore_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = uncore_io_mem_axi_0_r_ready;
  assign io_mmio_axi_0_aw_valid = uncore_io_mmio_axi_0_aw_valid;
  assign io_mmio_axi_0_aw_bits_addr = uncore_io_mmio_axi_0_aw_bits_addr;
  assign io_mmio_axi_0_aw_bits_len = uncore_io_mmio_axi_0_aw_bits_len;
  assign io_mmio_axi_0_aw_bits_size = uncore_io_mmio_axi_0_aw_bits_size;
  assign io_mmio_axi_0_aw_bits_burst = uncore_io_mmio_axi_0_aw_bits_burst;
  assign io_mmio_axi_0_aw_bits_lock = uncore_io_mmio_axi_0_aw_bits_lock;
  assign io_mmio_axi_0_aw_bits_cache = uncore_io_mmio_axi_0_aw_bits_cache;
  assign io_mmio_axi_0_aw_bits_prot = uncore_io_mmio_axi_0_aw_bits_prot;
  assign io_mmio_axi_0_aw_bits_qos = uncore_io_mmio_axi_0_aw_bits_qos;
  assign io_mmio_axi_0_aw_bits_region = uncore_io_mmio_axi_0_aw_bits_region;
  assign io_mmio_axi_0_aw_bits_id = uncore_io_mmio_axi_0_aw_bits_id;
  assign io_mmio_axi_0_aw_bits_user = uncore_io_mmio_axi_0_aw_bits_user;
  assign io_mmio_axi_0_w_valid = uncore_io_mmio_axi_0_w_valid;
  assign io_mmio_axi_0_w_bits_data = uncore_io_mmio_axi_0_w_bits_data;
  assign io_mmio_axi_0_w_bits_last = uncore_io_mmio_axi_0_w_bits_last;
  assign io_mmio_axi_0_w_bits_id = uncore_io_mmio_axi_0_w_bits_id;
  assign io_mmio_axi_0_w_bits_strb = uncore_io_mmio_axi_0_w_bits_strb;
  assign io_mmio_axi_0_w_bits_user = uncore_io_mmio_axi_0_w_bits_user;
  assign io_mmio_axi_0_b_ready = uncore_io_mmio_axi_0_b_ready;
  assign io_mmio_axi_0_ar_valid = uncore_io_mmio_axi_0_ar_valid;
  assign io_mmio_axi_0_ar_bits_addr = uncore_io_mmio_axi_0_ar_bits_addr;
  assign io_mmio_axi_0_ar_bits_len = uncore_io_mmio_axi_0_ar_bits_len;
  assign io_mmio_axi_0_ar_bits_size = uncore_io_mmio_axi_0_ar_bits_size;
  assign io_mmio_axi_0_ar_bits_burst = uncore_io_mmio_axi_0_ar_bits_burst;
  assign io_mmio_axi_0_ar_bits_lock = uncore_io_mmio_axi_0_ar_bits_lock;
  assign io_mmio_axi_0_ar_bits_cache = uncore_io_mmio_axi_0_ar_bits_cache;
  assign io_mmio_axi_0_ar_bits_prot = uncore_io_mmio_axi_0_ar_bits_prot;
  assign io_mmio_axi_0_ar_bits_qos = uncore_io_mmio_axi_0_ar_bits_qos;
  assign io_mmio_axi_0_ar_bits_region = uncore_io_mmio_axi_0_ar_bits_region;
  assign io_mmio_axi_0_ar_bits_id = uncore_io_mmio_axi_0_ar_bits_id;
  assign io_mmio_axi_0_ar_bits_user = uncore_io_mmio_axi_0_ar_bits_user;
  assign io_mmio_axi_0_r_ready = uncore_io_mmio_axi_0_r_ready;
  assign io_debug_req_ready = uncore_io_debugBus_req_ready;
  assign io_debug_resp_valid = uncore_io_debugBus_resp_valid;
  assign io_debug_resp_bits_resp = uncore_io_debugBus_resp_bits_resp;
  assign io_debug_resp_bits_data = uncore_io_debugBus_resp_bits_data;
  assign tileResets_0 = uncore_io_prci_0_reset;
  assign RocketTile_1_clk = clk;
  assign RocketTile_1_reset = tileResets_0;
  assign RocketTile_1_io_cached_0_acquire_ready = uncore_io_tiles_cached_0_acquire_ready;
  assign RocketTile_1_io_cached_0_probe_valid = uncore_io_tiles_cached_0_probe_valid;
  assign RocketTile_1_io_cached_0_probe_bits_addr_block = uncore_io_tiles_cached_0_probe_bits_addr_block;
  assign RocketTile_1_io_cached_0_probe_bits_p_type = uncore_io_tiles_cached_0_probe_bits_p_type;
  assign RocketTile_1_io_cached_0_release_ready = uncore_io_tiles_cached_0_release_ready;
  assign RocketTile_1_io_cached_0_grant_valid = uncore_io_tiles_cached_0_grant_valid;
  assign RocketTile_1_io_cached_0_grant_bits_addr_beat = uncore_io_tiles_cached_0_grant_bits_addr_beat;
  assign RocketTile_1_io_cached_0_grant_bits_client_xact_id = uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  assign RocketTile_1_io_cached_0_grant_bits_manager_xact_id = uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign RocketTile_1_io_cached_0_grant_bits_is_builtin_type = uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign RocketTile_1_io_cached_0_grant_bits_g_type = uncore_io_tiles_cached_0_grant_bits_g_type;
  assign RocketTile_1_io_cached_0_grant_bits_data = uncore_io_tiles_cached_0_grant_bits_data;
  assign RocketTile_1_io_cached_0_grant_bits_manager_id = uncore_io_tiles_cached_0_grant_bits_manager_id;
  assign RocketTile_1_io_cached_0_finish_ready = uncore_io_tiles_cached_0_finish_ready;
  assign RocketTile_1_io_uncached_0_acquire_ready = uncore_io_tiles_uncached_0_acquire_ready;
  assign RocketTile_1_io_uncached_0_grant_valid = uncore_io_tiles_uncached_0_grant_valid;
  assign RocketTile_1_io_uncached_0_grant_bits_addr_beat = uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  assign RocketTile_1_io_uncached_0_grant_bits_client_xact_id = uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign RocketTile_1_io_uncached_0_grant_bits_manager_xact_id = uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign RocketTile_1_io_uncached_0_grant_bits_is_builtin_type = uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign RocketTile_1_io_uncached_0_grant_bits_g_type = uncore_io_tiles_uncached_0_grant_bits_g_type;
  assign RocketTile_1_io_uncached_0_grant_bits_data = uncore_io_tiles_uncached_0_grant_bits_data;
  assign RocketTile_1_io_prci_reset = uncore_io_prci_0_reset;
  assign RocketTile_1_io_prci_id = uncore_io_prci_0_id;
  assign RocketTile_1_io_prci_interrupts_meip = uncore_io_prci_0_interrupts_meip;
  assign RocketTile_1_io_prci_interrupts_seip = uncore_io_prci_0_interrupts_seip;
  assign RocketTile_1_io_prci_interrupts_debug = uncore_io_prci_0_interrupts_debug;
  assign RocketTile_1_io_prci_interrupts_mtip = uncore_io_prci_0_interrupts_mtip;
  assign RocketTile_1_io_prci_interrupts_msip = uncore_io_prci_0_interrupts_msip;
  assign uncore_clk = clk;
  assign uncore_reset = reset;
  assign uncore_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign uncore_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign uncore_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign uncore_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign uncore_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign uncore_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign uncore_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign uncore_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign uncore_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign uncore_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign uncore_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign uncore_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign uncore_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign uncore_io_tiles_cached_0_acquire_valid = RocketTile_1_io_cached_0_acquire_valid;
  assign uncore_io_tiles_cached_0_acquire_bits_addr_block = RocketTile_1_io_cached_0_acquire_bits_addr_block;
  assign uncore_io_tiles_cached_0_acquire_bits_client_xact_id = RocketTile_1_io_cached_0_acquire_bits_client_xact_id;
  assign uncore_io_tiles_cached_0_acquire_bits_addr_beat = RocketTile_1_io_cached_0_acquire_bits_addr_beat;
  assign uncore_io_tiles_cached_0_acquire_bits_is_builtin_type = RocketTile_1_io_cached_0_acquire_bits_is_builtin_type;
  assign uncore_io_tiles_cached_0_acquire_bits_a_type = RocketTile_1_io_cached_0_acquire_bits_a_type;
  assign uncore_io_tiles_cached_0_acquire_bits_union = RocketTile_1_io_cached_0_acquire_bits_union;
  assign uncore_io_tiles_cached_0_acquire_bits_data = RocketTile_1_io_cached_0_acquire_bits_data;
  assign uncore_io_tiles_cached_0_probe_ready = RocketTile_1_io_cached_0_probe_ready;
  assign uncore_io_tiles_cached_0_release_valid = RocketTile_1_io_cached_0_release_valid;
  assign uncore_io_tiles_cached_0_release_bits_addr_beat = RocketTile_1_io_cached_0_release_bits_addr_beat;
  assign uncore_io_tiles_cached_0_release_bits_addr_block = RocketTile_1_io_cached_0_release_bits_addr_block;
  assign uncore_io_tiles_cached_0_release_bits_client_xact_id = RocketTile_1_io_cached_0_release_bits_client_xact_id;
  assign uncore_io_tiles_cached_0_release_bits_voluntary = RocketTile_1_io_cached_0_release_bits_voluntary;
  assign uncore_io_tiles_cached_0_release_bits_r_type = RocketTile_1_io_cached_0_release_bits_r_type;
  assign uncore_io_tiles_cached_0_release_bits_data = RocketTile_1_io_cached_0_release_bits_data;
  assign uncore_io_tiles_cached_0_grant_ready = RocketTile_1_io_cached_0_grant_ready;
  assign uncore_io_tiles_cached_0_finish_valid = RocketTile_1_io_cached_0_finish_valid;
  assign uncore_io_tiles_cached_0_finish_bits_manager_xact_id = RocketTile_1_io_cached_0_finish_bits_manager_xact_id;
  assign uncore_io_tiles_cached_0_finish_bits_manager_id = RocketTile_1_io_cached_0_finish_bits_manager_id;
  assign uncore_io_tiles_uncached_0_acquire_valid = RocketTile_1_io_uncached_0_acquire_valid;
  assign uncore_io_tiles_uncached_0_acquire_bits_addr_block = RocketTile_1_io_uncached_0_acquire_bits_addr_block;
  assign uncore_io_tiles_uncached_0_acquire_bits_client_xact_id = RocketTile_1_io_uncached_0_acquire_bits_client_xact_id;
  assign uncore_io_tiles_uncached_0_acquire_bits_addr_beat = RocketTile_1_io_uncached_0_acquire_bits_addr_beat;
  assign uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type = RocketTile_1_io_uncached_0_acquire_bits_is_builtin_type;
  assign uncore_io_tiles_uncached_0_acquire_bits_a_type = RocketTile_1_io_uncached_0_acquire_bits_a_type;
  assign uncore_io_tiles_uncached_0_acquire_bits_union = RocketTile_1_io_uncached_0_acquire_bits_union;
  assign uncore_io_tiles_uncached_0_acquire_bits_data = RocketTile_1_io_uncached_0_acquire_bits_data;
  assign uncore_io_tiles_uncached_0_grant_ready = RocketTile_1_io_uncached_0_grant_ready;
  assign uncore_io_mmio_axi_0_aw_ready = io_mmio_axi_0_aw_ready;
  assign uncore_io_mmio_axi_0_w_ready = io_mmio_axi_0_w_ready;
  assign uncore_io_mmio_axi_0_b_valid = io_mmio_axi_0_b_valid;
  assign uncore_io_mmio_axi_0_b_bits_resp = io_mmio_axi_0_b_bits_resp;
  assign uncore_io_mmio_axi_0_b_bits_id = io_mmio_axi_0_b_bits_id;
  assign uncore_io_mmio_axi_0_b_bits_user = io_mmio_axi_0_b_bits_user;
  assign uncore_io_mmio_axi_0_ar_ready = io_mmio_axi_0_ar_ready;
  assign uncore_io_mmio_axi_0_r_valid = io_mmio_axi_0_r_valid;
  assign uncore_io_mmio_axi_0_r_bits_resp = io_mmio_axi_0_r_bits_resp;
  assign uncore_io_mmio_axi_0_r_bits_data = io_mmio_axi_0_r_bits_data;
  assign uncore_io_mmio_axi_0_r_bits_last = io_mmio_axi_0_r_bits_last;
  assign uncore_io_mmio_axi_0_r_bits_id = io_mmio_axi_0_r_bits_id;
  assign uncore_io_mmio_axi_0_r_bits_user = io_mmio_axi_0_r_bits_user;
  assign uncore_io_interrupts_0 = io_interrupts_0;
  assign uncore_io_interrupts_1 = io_interrupts_1;
  assign uncore_io_debugBus_req_valid = io_debug_req_valid;
  assign uncore_io_debugBus_req_bits_addr = io_debug_req_bits_addr;
  assign uncore_io_debugBus_req_bits_op = io_debug_req_bits_op;
  assign uncore_io_debugBus_req_bits_data = io_debug_req_bits_data;
  assign uncore_io_debugBus_resp_ready = io_debug_resp_ready;
endmodule
